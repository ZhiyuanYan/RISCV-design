module top(input rst,
	input clk,
	input [34:0] i44,
	input [4:0] i41,
	input [4:0] i40,
	input [31:0] i39,
	input [34:0] i42,
	input [31:0] i38,
	input [3:0] i36,
	input [31:0] i35,
	input [36:0] i43,
	input [15:0] i34,
	input [15:0] i33,
	input [31:0] i32,
	input [23:0] i31,
	input [31:0] i11,
	input [31:0] i18,
	input [7:0] i48,
	input [31:0] i10,
	input [31:0] i37,
	input [0:0] i9,
	input [2:0] i15,
	input [0:0] i8,
	input [7:0] i47,
	input [0:0] i7,
	input [1:0] i23,
	input [0:0] i21,
	input [31:0] i6,
	input [0:0] i5,
	input [31:0] i45,
	input [31:0] i27,
	input [0:0] i4,
	input [31:0] i26,
	input [0:0] i17,
	input [2:0] i16,
	input [0:0] i3,
	input [0:0] i2,
	input [23:0] i30,
	input [0:0] i1,
	input [0:0] i12,
	input [0:0] i0,
	input [0:0] i13,
	input [31:0] i14,
	input [0:0] i19,
	input [31:0] i20,
	input [31:0] i46,
	input [23:0] i29,
	input [23:0] i28,
	input [1:0] i22,
	input [1:0] i24,
	input [31:0] i25,
	output [31:0] o11,
	output [0:0] o10,
	output [3:0] o9,
	output [31:0] o8,
	output [0:0] o7,
	output [0:0] o12,
	output [2:0] o4,
	output [31:0] o3,
	output [0:0] o2,
	output [0:0] o6,
	output [0:0] o5,
	output [2:0] o1,
	output [31:0] o0
);

	// states
	reg [31:0] s18;
	reg [31:0] s19;
	reg [1:0] s22;
	reg [31:0] s31;
	reg [3:0] s49;
	reg [0:0] s55;
	reg [31:0] s107;
	reg [3:0] s109;
	reg [31:0] s118;
	reg [0:0] s121;
	reg [0:0] s123;
	reg [11:0] s127;
	reg [0:0] s152;
	reg [0:0] s180;
	reg [1:0] s235;
	reg [0:0] s239;
	reg [0:0] s297;
	reg [31:0] s302;
	reg [31:0] s305;
	reg [15:0] s404;
	reg [15:0] s409;
	reg [31:0] s415;
	reg [31:0] s416;
	reg [31:0] s417;
	reg [31:0] s418;
	reg [31:0] s419;
	reg [31:0] s420;
	reg [31:0] s421;
	reg [31:0] s422;
	reg [31:0] s437;
	reg [31:0] s438;
	reg [31:0] s439;
	reg [31:0] s440;
	reg [31:0] s441;
	reg [31:0] s442;
	reg [31:0] s443;
	reg [31:0] s444;
	reg [31:0] s453;
	reg [31:0] s454;
	reg [31:0] s455;
	reg [31:0] s456;
	reg [31:0] s457;
	reg [31:0] s458;
	reg [31:0] s459;
	reg [31:0] s460;
	reg [31:0] s468;
	reg [31:0] s469;
	reg [31:0] s470;
	reg [31:0] s471;
	reg [31:0] s472;
	reg [31:0] s473;
	reg [31:0] s474;
	reg [31:0] s475;
	reg [31:0] s762;
	reg [31:0] s769;
	reg [0:0] s772;
	reg [6:0] s792;
	reg [6:0] s797;
	reg [31:0] s813;
	reg [31:0] s815;
	reg [1:0] s885;
	reg [0:0] s896;
	reg [0:0] s898;
	reg [0:0] s900;
	reg [32:0] s960;
	reg [31:0] s984;
	reg [63:0] s1004;
	reg [63:0] s1007;
	reg [63:0] s1009;
	reg [63:0] s1011;
	reg [63:0] s1043;
	reg [31:0] s1066;
	reg [31:0] s1069;
	reg [1:0] s1127;
	reg [4:0] s1134;
	reg [34:0] s1160;
	reg [16:0] s1191;
	reg [1:0] s1201;
	reg [4:0] s1207;
	reg [36:0] s1234;
	reg [17:0] s1254;
	reg [1:0] s1264;
	reg [4:0] s1270;
	reg [34:0] s1294;
	reg [16:0] s1305;
	reg [63:0] s1467;
	reg [31:0] s1490;
	reg [31:0] s1491;
	reg [6:0] s1492;
	reg [31:0] s1496;
	reg [31:0] s1497;
	reg [31:0] s1501;
	reg [31:0] s1502;
	reg [31:0] s1504;
	reg [31:0] s1505;
	reg [31:0] s1510;
	reg [31:0] s1511;
	reg [31:0] s1513;
	reg [31:0] s1514;
	reg [31:0] s1517;
	reg [31:0] s1518;
	reg [31:0] s1520;
	reg [31:0] s1521;
	reg [31:0] s1527;
	reg [31:0] s1528;
	reg [31:0] s1530;
	reg [31:0] s1531;
	reg [31:0] s1534;
	reg [31:0] s1535;
	reg [31:0] s1537;
	reg [31:0] s1538;
	reg [31:0] s1542;
	reg [31:0] s1543;
	reg [31:0] s1545;
	reg [31:0] s1546;
	reg [31:0] s1549;
	reg [31:0] s1550;
	reg [31:0] s1552;
	reg [31:0] s1553;
	reg [31:0] s1560;
	reg [31:0] s1561;
	reg [31:0] s1563;
	reg [31:0] s1564;
	reg [31:0] s1567;
	reg [31:0] s1568;
	reg [31:0] s1570;
	reg [31:0] s1571;
	reg [31:0] s1575;
	reg [31:0] s1576;
	reg [31:0] s1578;
	reg [31:0] s1579;
	reg [31:0] s1582;
	reg [31:0] s1583;
	reg [31:0] s1585;
	reg [31:0] s1586;
	reg [31:0] s1591;
	reg [31:0] s1592;
	reg [31:0] s1594;
	reg [31:0] s1595;
	reg [31:0] s1598;
	reg [31:0] s1599;
	reg [31:0] s1601;
	reg [31:0] s1602;
	reg [31:0] s1606;
	reg [31:0] s1607;
	reg [31:0] s1609;
	reg [31:0] s1610;
	reg [31:0] s1613;
	reg [31:0] s1614;
	reg [31:0] s1616;
	reg [31:0] s1617;
	reg [31:0] s1625;
	reg [31:0] s1626;
	reg [31:0] s1628;
	reg [31:0] s1629;
	reg [31:0] s1632;
	reg [31:0] s1633;
	reg [31:0] s1635;
	reg [31:0] s1636;
	reg [31:0] s1640;
	reg [31:0] s1641;
	reg [31:0] s1643;
	reg [31:0] s1644;
	reg [31:0] s1647;
	reg [31:0] s1648;
	reg [31:0] s1650;
	reg [31:0] s1651;
	reg [31:0] s1656;
	reg [31:0] s1657;
	reg [31:0] s1659;
	reg [31:0] s1660;
	reg [31:0] s1663;
	reg [31:0] s1664;
	reg [31:0] s1666;
	reg [31:0] s1667;
	reg [31:0] s1671;
	reg [31:0] s1672;
	reg [31:0] s1674;
	reg [31:0] s1675;
	reg [31:0] s1678;
	reg [31:0] s1679;
	reg [31:0] s1681;
	reg [31:0] s1682;
	reg [31:0] s1688;
	reg [31:0] s1689;
	reg [31:0] s1691;
	reg [31:0] s1692;
	reg [31:0] s1695;
	reg [31:0] s1696;
	reg [31:0] s1698;
	reg [31:0] s1699;
	reg [31:0] s1703;
	reg [31:0] s1704;
	reg [31:0] s1706;
	reg [31:0] s1707;
	reg [31:0] s1710;
	reg [31:0] s1711;
	reg [31:0] s1713;
	reg [31:0] s1714;
	reg [31:0] s1719;
	reg [31:0] s1720;
	reg [31:0] s1722;
	reg [31:0] s1723;
	reg [31:0] s1726;
	reg [31:0] s1727;
	reg [31:0] s1729;
	reg [31:0] s1730;
	reg [31:0] s1734;
	reg [31:0] s1735;
	reg [31:0] s1737;
	reg [31:0] s1738;
	reg [31:0] s1741;
	reg [31:0] s1742;
	reg [31:0] s1744;
	reg [31:0] s1745;
	reg [31:0] s1754;
	reg [31:0] s1755;
	reg [31:0] s1757;
	reg [31:0] s1758;
	reg [31:0] s1761;
	reg [31:0] s1762;
	reg [31:0] s1764;
	reg [31:0] s1765;
	reg [31:0] s1769;
	reg [31:0] s1770;
	reg [31:0] s1772;
	reg [31:0] s1773;
	reg [31:0] s1776;
	reg [31:0] s1777;
	reg [31:0] s1779;
	reg [31:0] s1780;
	reg [31:0] s1785;
	reg [31:0] s1786;
	reg [31:0] s1788;
	reg [31:0] s1789;
	reg [31:0] s1792;
	reg [31:0] s1793;
	reg [31:0] s1795;
	reg [31:0] s1796;
	reg [31:0] s1800;
	reg [31:0] s1801;
	reg [31:0] s1803;
	reg [31:0] s1804;
	reg [31:0] s1807;
	reg [31:0] s1808;
	reg [31:0] s1810;
	reg [31:0] s1811;
	reg [31:0] s1817;
	reg [31:0] s1818;
	reg [31:0] s1820;
	reg [31:0] s1821;
	reg [31:0] s1824;
	reg [31:0] s1825;
	reg [31:0] s1827;
	reg [31:0] s1828;
	reg [31:0] s1832;
	reg [31:0] s1833;
	reg [31:0] s1835;
	reg [31:0] s1836;
	reg [31:0] s1839;
	reg [31:0] s1840;
	reg [31:0] s1842;
	reg [31:0] s1843;
	reg [31:0] s1848;
	reg [31:0] s1849;
	reg [31:0] s1851;
	reg [31:0] s1852;
	reg [31:0] s1855;
	reg [31:0] s1856;
	reg [31:0] s1858;
	reg [31:0] s1859;
	reg [31:0] s1863;
	reg [31:0] s1864;
	reg [31:0] s1866;
	reg [31:0] s1867;
	reg [31:0] s1870;
	reg [31:0] s1871;
	reg [31:0] s1873;
	reg [31:0] s1874;
	reg [31:0] s1881;
	reg [31:0] s1882;
	reg [31:0] s1884;
	reg [31:0] s1885;
	reg [31:0] s1888;
	reg [31:0] s1889;
	reg [31:0] s1891;
	reg [31:0] s1892;
	reg [31:0] s1896;
	reg [31:0] s1897;
	reg [31:0] s1899;
	reg [31:0] s1900;
	reg [31:0] s1903;
	reg [31:0] s1904;
	reg [31:0] s1906;
	reg [31:0] s1907;
	reg [31:0] s1912;
	reg [31:0] s1913;
	reg [31:0] s1915;
	reg [31:0] s1916;
	reg [31:0] s1919;
	reg [31:0] s1920;
	reg [31:0] s1922;
	reg [31:0] s1923;
	reg [31:0] s1927;
	reg [31:0] s1928;
	reg [31:0] s1930;
	reg [31:0] s1931;
	reg [31:0] s1934;
	reg [31:0] s1935;
	reg [31:0] s1937;
	reg [31:0] s1938;
	reg [31:0] s1944;
	reg [31:0] s1945;
	reg [31:0] s1947;
	reg [31:0] s1948;
	reg [31:0] s1951;
	reg [31:0] s1952;
	reg [31:0] s1954;
	reg [31:0] s1955;
	reg [31:0] s1959;
	reg [31:0] s1960;
	reg [31:0] s1962;
	reg [31:0] s1963;
	reg [31:0] s1966;
	reg [31:0] s1967;
	reg [31:0] s1969;
	reg [31:0] s1970;
	reg [31:0] s1975;
	reg [31:0] s1976;
	reg [31:0] s1978;
	reg [31:0] s1979;
	reg [31:0] s1982;
	reg [31:0] s1983;
	reg [31:0] s1985;
	reg [31:0] s1986;
	reg [31:0] s1990;
	reg [31:0] s1991;
	reg [31:0] s1993;
	reg [31:0] s1994;
	reg [31:0] s1997;
	reg [31:0] s1998;
	reg [31:0] s2000;
	reg [31:0] s2001;
	reg [31:0] s2596;
	reg [31:0] s2597;
	reg [0:0] s2600;
	reg [0:0] s2601;
	reg [31:0] s2604;
	reg [31:0] s2606;
	reg [0:0] s2609;
	reg [0:0] s2611;
	reg [0:0] s2612;
	reg [0:0] s2615;
	reg [31:0] s2617;
	reg [31:0] s2618;
	reg [31:0] s2624;
	reg [31:0] s2626;
	reg [31:0] s2632;
	reg [0:0] s2700;
	reg [0:0] s2702;
	reg [31:0] s2705;
	reg [31:0] s2729;
	reg [3:0] s2760;
	reg [31:0] s2971;
	reg [31:0] s2991;
	reg [0:0] s2995;
	reg [4:0] s2997;
	reg [31:0] s2999;
	reg [31:0] s3000;
	reg [31:0] s3001;
	reg [31:0] s3006;
	reg [31:0] s3011;
	reg [31:0] s3038;
	reg [31:0] s3040;
	reg [31:0] s3045;
	reg [31:0] s3047;

	// wires
	wire [31:0] w20;
	wire [0:0] w23;
	wire [1:0] w24;
	wire [0:0] w25;
	wire [0:0] w26;
	wire [0:0] w27;
	wire [1:0] w28;
	wire [0:0] w29;
	wire [31:0] w30;
	wire [1:0] w32;
	wire [0:0] w33;
	wire [1:0] w34;
	wire [0:0] w35;
	wire [1:0] w36;
	wire [0:0] w37;
	wire [31:0] w38;
	wire [2:0] w42;
	wire [2:0] w43;
	wire [2:0] w44;
	wire [2:0] w45;
	wire [0:0] w47;
	wire [3:0] w50;
	wire [0:0] w51;
	wire [0:0] w52;
	wire [0:0] w53;
	wire [0:0] w54;
	wire [0:0] w56;
	wire [0:0] w57;
	wire [0:0] w58;
	wire [0:0] w59;
	wire [0:0] w60;
	wire [0:0] w61;
	wire [1:0] w65;
	wire [2:0] w66;
	wire [3:0] w67;
	wire [0:0] w68;
	wire [2:0] w69;
	wire [2:0] w71;
	wire [3:0] w72;
	wire [0:0] w73;
	wire [2:0] w74;
	wire [3:0] w75;
	wire [0:0] w76;
	wire [1:0] w77;
	wire [0:0] w78;
	wire [0:0] w79;
	wire [0:0] w80;
	wire [0:0] w81;
	wire [0:0] w82;
	wire [0:0] w83;
	wire [0:0] w84;
	wire [3:0] w86;
	wire [0:0] w87;
	wire [2:0] w88;
	wire [3:0] w89;
	wire [0:0] w90;
	wire [1:0] w91;
	wire [2:0] w92;
	wire [3:0] w93;
	wire [0:0] w94;
	wire [0:0] w95;
	wire [0:0] w96;
	wire [0:0] w97;
	wire [3:0] w99;
	wire [0:0] w100;
	wire [1:0] w101;
	wire [0:0] w102;
	wire [0:0] w103;
	wire [0:0] w104;
	wire [0:0] w105;
	wire [1:0] w111;
	wire [0:0] w112;
	wire [0:0] w113;
	wire [0:0] w114;
	wire [0:0] w115;
	wire [31:0] w117;
	wire [0:0] w125;
	wire [6:0] w129;
	wire [11:0] w130;
	wire [0:0] w131;
	wire [6:0] w132;
	wire [11:0] w133;
	wire [0:0] w134;
	wire [5:0] w136;
	wire [11:0] w137;
	wire [0:0] w138;
	wire [4:0] w140;
	wire [11:0] w141;
	wire [0:0] w142;
	wire [6:0] w143;
	wire [11:0] w144;
	wire [0:0] w145;
	wire [1:0] w146;
	wire [2:0] w147;
	wire [3:0] w148;
	wire [4:0] w149;
	wire [0:0] w150;
	wire [0:0] w151;
	wire [10:0] w154;
	wire [11:0] w155;
	wire [0:0] w156;
	wire [11:0] w157;
	wire [0:0] w158;
	wire [7:0] w160;
	wire [11:0] w161;
	wire [0:0] w162;
	wire [7:0] w163;
	wire [11:0] w164;
	wire [0:0] w165;
	wire [9:0] w167;
	wire [11:0] w168;
	wire [0:0] w169;
	wire [9:0] w170;
	wire [11:0] w171;
	wire [0:0] w172;
	wire [1:0] w173;
	wire [2:0] w174;
	wire [3:0] w175;
	wire [4:0] w176;
	wire [5:0] w177;
	wire [0:0] w178;
	wire [0:0] w179;
	wire [5:0] w181;
	wire [11:0] w182;
	wire [0:0] w183;
	wire [4:0] w184;
	wire [11:0] w185;
	wire [0:0] w186;
	wire [8:0] w188;
	wire [11:0] w189;
	wire [0:0] w190;
	wire [8:0] w191;
	wire [11:0] w192;
	wire [0:0] w193;
	wire [8:0] w194;
	wire [11:0] w195;
	wire [0:0] w196;
	wire [8:0] w197;
	wire [11:0] w198;
	wire [0:0] w199;
	wire [9:0] w200;
	wire [11:0] w201;
	wire [0:0] w202;
	wire [9:0] w203;
	wire [11:0] w204;
	wire [0:0] w205;
	wire [9:0] w206;
	wire [11:0] w207;
	wire [0:0] w208;
	wire [9:0] w209;
	wire [11:0] w210;
	wire [0:0] w211;
	wire [9:0] w212;
	wire [11:0] w213;
	wire [0:0] w214;
	wire [9:0] w215;
	wire [11:0] w216;
	wire [0:0] w217;
	wire [11:0] w218;
	wire [0:0] w219;
	wire [1:0] w220;
	wire [2:0] w221;
	wire [3:0] w222;
	wire [4:0] w223;
	wire [5:0] w224;
	wire [6:0] w225;
	wire [7:0] w226;
	wire [8:0] w227;
	wire [9:0] w228;
	wire [10:0] w229;
	wire [11:0] w230;
	wire [12:0] w232;
	wire [0:0] w233;
	wire [0:0] w234;
	wire [0:0] w236;
	wire [0:0] w237;
	wire [0:0] w238;
	wire [0:0] w240;
	wire [0:0] w242;
	wire [0:0] w243;
	wire [0:0] w244;
	wire [0:0] w245;
	wire [0:0] w246;
	wire [0:0] w247;
	wire [0:0] w248;
	wire [0:0] w249;
	wire [0:0] w250;
	wire [0:0] w251;
	wire [1:0] w252;
	wire [2:0] w253;
	wire [0:0] w254;
	wire [0:0] w255;
	wire [0:0] w256;
	wire [0:0] w257;
	wire [0:0] w258;
	wire [0:0] w259;
	wire [0:0] w260;
	wire [0:0] w261;
	wire [0:0] w262;
	wire [0:0] w263;
	wire [0:0] w264;
	wire [0:0] w265;
	wire [0:0] w266;
	wire [0:0] w267;
	wire [0:0] w268;
	wire [0:0] w269;
	wire [0:0] w270;
	wire [0:0] w271;
	wire [0:0] w272;
	wire [0:0] w273;
	wire [0:0] w274;
	wire [0:0] w275;
	wire [0:0] w276;
	wire [0:0] w277;
	wire [0:0] w278;
	wire [0:0] w279;
	wire [0:0] w280;
	wire [0:0] w281;
	wire [0:0] w282;
	wire [0:0] w283;
	wire [0:0] w284;
	wire [0:0] w285;
	wire [0:0] w286;
	wire [0:0] w287;
	wire [0:0] w288;
	wire [0:0] w289;
	wire [0:0] w290;
	wire [0:0] w291;
	wire [0:0] w292;
	wire [0:0] w293;
	wire [0:0] w294;
	wire [0:0] w295;
	wire [0:0] w296;
	wire [0:0] w298;
	wire [0:0] w299;
	wire [0:0] w300;
	wire [4:0] w301;
	wire [31:0] w303;
	wire [31:0] w304;
	wire [4:0] w307;
	wire [2:0] w308;
	wire [0:0] w309;
	wire [4:0] w310;
	wire [6:0] w311;
	wire [4:0] w312;
	wire [6:0] w313;
	wire [0:0] w314;
	wire [4:0] w315;
	wire [0:0] w316;
	wire [4:0] w317;
	wire [0:0] w318;
	wire [0:0] w319;
	wire [4:0] w320;
	wire [0:0] w321;
	wire [4:0] w322;
	wire [4:0] w323;
	wire [0:0] w324;
	wire [5:0] w325;
	wire [0:0] w326;
	wire [0:0] w327;
	wire [6:0] w328;
	wire [6:0] w329;
	wire [0:0] w330;
	wire [0:0] w331;
	wire [0:0] w332;
	wire [0:0] w333;
	wire [0:0] w334;
	wire [4:0] w335;
	wire [6:0] w336;
	wire [0:0] w337;
	wire [4:0] w338;
	wire [6:0] w339;
	wire [0:0] w340;
	wire [4:0] w341;
	wire [1:0] w342;
	wire [0:0] w343;
	wire [0:0] w344;
	wire [4:0] w345;
	wire [5:0] w346;
	wire [6:0] w347;
	wire [0:0] w348;
	wire [4:0] w349;
	wire [1:0] w350;
	wire [0:0] w351;
	wire [0:0] w352;
	wire [4:0] w353;
	wire [6:0] w354;
	wire [0:0] w355;
	wire [4:0] w356;
	wire [0:0] w357;
	wire [0:0] w358;
	wire [0:0] w359;
	wire [4:0] w360;
	wire [6:0] w361;
	wire [0:0] w362;
	wire [4:0] w363;
	wire [4:0] w364;
	wire [0:0] w365;
	wire [4:0] w366;
	wire [4:0] w367;
	wire [0:0] w368;
	wire [6:0] w369;
	wire [0:0] w370;
	wire [6:0] w371;
	wire [0:0] w372;
	wire [1:0] w373;
	wire [2:0] w374;
	wire [0:0] w375;
	wire [4:0] w376;
	wire [4:0] w377;
	wire [4:0] w378;
	wire [4:0] w379;
	wire [4:0] w380;
	wire [4:0] w381;
	wire [4:0] w382;
	wire [4:0] w383;
	wire [4:0] w384;
	wire [1:0] w385;
	wire [2:0] w386;
	wire [3:0] w387;
	wire [0:0] w388;
	wire [4:0] w389;
	wire [4:0] w390;
	wire [4:0] w391;
	wire [4:0] w392;
	wire [4:0] w393;
	wire [4:0] w394;
	wire [4:0] w395;
	wire [4:0] w396;
	wire [4:0] w397;
	wire [4:0] w398;
	wire [0:0] w399;
	wire [0:0] w400;
	wire [0:0] w401;
	wire [15:0] w403;
	wire [0:0] w406;
	wire [0:0] w407;
	wire [0:0] w408;
	wire [0:0] w411;
	wire [0:0] w412;
	wire [0:0] w413;
	wire [0:0] w414;
	wire [63:0] w424;
	wire [95:0] w426;
	wire [127:0] w428;
	wire [159:0] w430;
	wire [191:0] w432;
	wire [223:0] w434;
	wire [255:0] w436;
	wire [63:0] w445;
	wire [95:0] w446;
	wire [127:0] w447;
	wire [159:0] w448;
	wire [191:0] w449;
	wire [223:0] w450;
	wire [255:0] w451;
	wire [255:0] w452;
	wire [63:0] w461;
	wire [95:0] w462;
	wire [127:0] w463;
	wire [159:0] w464;
	wire [191:0] w465;
	wire [223:0] w466;
	wire [255:0] w467;
	wire [63:0] w476;
	wire [95:0] w477;
	wire [127:0] w478;
	wire [159:0] w479;
	wire [191:0] w480;
	wire [223:0] w481;
	wire [255:0] w482;
	wire [255:0] w483;
	wire [255:0] w484;
	wire [31:0] w485;
	wire [255:0] w486;
	wire [255:0] w487;
	wire [255:0] w488;
	wire [31:0] w489;
	wire [0:0] w490;
	wire [31:0] w491;
	wire [31:0] w492;
	wire [0:0] w493;
	wire [0:0] w494;
	wire [31:0] w495;
	wire [31:0] w496;
	wire [0:0] w497;
	wire [0:0] w498;
	wire [31:0] w499;
	wire [31:0] w500;
	wire [0:0] w501;
	wire [0:0] w502;
	wire [31:0] w503;
	wire [31:0] w504;
	wire [0:0] w505;
	wire [0:0] w506;
	wire [31:0] w507;
	wire [0:0] w508;
	wire [0:0] w509;
	wire [31:0] w510;
	wire [0:0] w511;
	wire [0:0] w512;
	wire [0:0] w513;
	wire [0:0] w514;
	wire [0:0] w515;
	wire [0:0] w516;
	wire [0:0] w517;
	wire [0:0] w518;
	wire [0:0] w519;
	wire [0:0] w520;
	wire [0:0] w521;
	wire [0:0] w522;
	wire [0:0] w523;
	wire [0:0] w524;
	wire [0:0] w525;
	wire [0:0] w526;
	wire [0:0] w527;
	wire [0:0] w528;
	wire [0:0] w529;
	wire [0:0] w530;
	wire [0:0] w531;
	wire [0:0] w532;
	wire [0:0] w533;
	wire [0:0] w535;
	wire [0:0] w536;
	wire [0:0] w537;
	wire [0:0] w538;
	wire [0:0] w539;
	wire [0:0] w540;
	wire [0:0] w541;
	wire [0:0] w542;
	wire [4:0] w543;
	wire [4:0] w544;
	wire [0:0] w545;
	wire [4:0] w546;
	wire [0:0] w547;
	wire [0:0] w548;
	wire [4:0] w549;
	wire [0:0] w550;
	wire [0:0] w551;
	wire [2:0] w552;
	wire [0:0] w553;
	wire [0:0] w554;
	wire [0:0] w555;
	wire [6:0] w556;
	wire [0:0] w557;
	wire [0:0] w558;
	wire [0:0] w559;
	wire [6:0] w560;
	wire [6:0] w561;
	wire [0:0] w562;
	wire [0:0] w563;
	wire [5:0] w564;
	wire [6:0] w565;
	wire [0:0] w566;
	wire [0:0] w567;
	wire [0:0] w568;
	wire [0:0] w569;
	wire [2:0] w570;
	wire [0:0] w571;
	wire [0:0] w572;
	wire [0:0] w573;
	wire [0:0] w574;
	wire [0:0] w575;
	wire [2:0] w576;
	wire [0:0] w577;
	wire [0:0] w578;
	wire [0:0] w579;
	wire [0:0] w580;
	wire [0:0] w581;
	wire [2:0] w582;
	wire [0:0] w583;
	wire [0:0] w584;
	wire [0:0] w585;
	wire [0:0] w586;
	wire [0:0] w587;
	wire [0:0] w588;
	wire [0:0] w589;
	wire [0:0] w590;
	wire [0:0] w591;
	wire [0:0] w592;
	wire [0:0] w593;
	wire [0:0] w594;
	wire [0:0] w595;
	wire [0:0] w596;
	wire [0:0] w597;
	wire [0:0] w598;
	wire [0:0] w599;
	wire [0:0] w600;
	wire [0:0] w601;
	wire [0:0] w602;
	wire [0:0] w603;
	wire [0:0] w604;
	wire [0:0] w605;
	wire [0:0] w606;
	wire [0:0] w607;
	wire [0:0] w608;
	wire [0:0] w609;
	wire [0:0] w610;
	wire [6:0] w611;
	wire [0:0] w612;
	wire [0:0] w613;
	wire [0:0] w614;
	wire [0:0] w615;
	wire [0:0] w616;
	wire [0:0] w617;
	wire [0:0] w618;
	wire [0:0] w619;
	wire [0:0] w620;
	wire [0:0] w621;
	wire [0:0] w622;
	wire [0:0] w623;
	wire [0:0] w624;
	wire [0:0] w625;
	wire [0:0] w626;
	wire [6:0] w627;
	wire [0:0] w628;
	wire [0:0] w629;
	wire [0:0] w630;
	wire [0:0] w631;
	wire [0:0] w632;
	wire [0:0] w633;
	wire [0:0] w634;
	wire [0:0] w635;
	wire [0:0] w636;
	wire [0:0] w637;
	wire [0:0] w638;
	wire [0:0] w639;
	wire [0:0] w640;
	wire [0:0] w641;
	wire [0:0] w642;
	wire [0:0] w643;
	wire [0:0] w644;
	wire [0:0] w645;
	wire [0:0] w646;
	wire [0:0] w647;
	wire [0:0] w648;
	wire [0:0] w649;
	wire [0:0] w650;
	wire [0:0] w651;
	wire [0:0] w652;
	wire [0:0] w653;
	wire [0:0] w654;
	wire [0:0] w655;
	wire [0:0] w656;
	wire [1:0] w657;
	wire [0:0] w658;
	wire [0:0] w659;
	wire [0:0] w660;
	wire [0:0] w661;
	wire [0:0] w662;
	wire [0:0] w663;
	wire [0:0] w664;
	wire [6:0] w665;
	wire [0:0] w666;
	wire [0:0] w667;
	wire [0:0] w668;
	wire [0:0] w669;
	wire [0:0] w670;
	wire [0:0] w671;
	wire [0:0] w672;
	wire [6:0] w673;
	wire [0:0] w674;
	wire [0:0] w675;
	wire [0:0] w676;
	wire [0:0] w677;
	wire [6:0] w678;
	wire [0:0] w679;
	wire [0:0] w680;
	wire [0:0] w681;
	wire [0:0] w682;
	wire [0:0] w684;
	wire [0:0] w685;
	wire [11:0] w687;
	wire [1:0] w688;
	wire [6:0] w689;
	wire [2:0] w690;
	wire [9:0] w691;
	wire [11:0] w692;
	wire [11:0] w693;
	wire [11:0] w694;
	wire [11:0] w695;
	wire [3:0] w696;
	wire [6:0] w697;
	wire [0:0] w698;
	wire [7:0] w699;
	wire [11:0] w700;
	wire [11:0] w701;
	wire [11:0] w702;
	wire [6:0] w703;
	wire [2:0] w704;
	wire [9:0] w705;
	wire [0:0] w706;
	wire [10:0] w707;
	wire [0:0] w708;
	wire [11:0] w709;
	wire [11:0] w710;
	wire [11:0] w711;
	wire [6:0] w712;
	wire [2:0] w713;
	wire [9:0] w714;
	wire [0:0] w715;
	wire [10:0] w716;
	wire [6:0] w717;
	wire [2:0] w718;
	wire [9:0] w719;
	wire [10:0] w720;
	wire [1:0] w721;
	wire [0:0] w722;
	wire [10:0] w723;
	wire [11:0] w724;
	wire [11:0] w725;
	wire [11:0] w726;
	wire [11:0] w727;
	wire [11:0] w728;
	wire [11:0] w729;
	wire [11:0] w730;
	wire [11:0] w731;
	wire [11:0] w732;
	wire [11:0] w733;
	wire [6:0] w734;
	wire [11:0] w735;
	wire [11:0] w736;
	wire [1:0] w737;
	wire [1:0] w738;
	wire [0:0] w739;
	wire [0:0] w740;
	wire [0:0] w741;
	wire [0:0] w742;
	wire [0:0] w743;
	wire [4:0] w744;
	wire [4:0] w745;
	wire [4:0] w746;
	wire [4:0] w747;
	wire [4:0] w748;
	wire [4:0] w749;
	wire [4:0] w750;
	wire [4:0] w751;
	wire [4:0] w752;
	wire [4:0] w753;
	wire [4:0] w754;
	wire [4:0] w755;
	wire [4:0] w756;
	wire [4:0] w757;
	wire [4:0] w758;
	wire [4:0] w759;
	wire [4:0] w760;
	wire [4:0] w761;
	wire [31:0] w763;
	wire [4:0] w764;
	wire [31:0] w765;
	wire [0:0] w766;
	wire [4:0] w767;
	wire [31:0] w770;
	wire [31:0] w771;
	wire [0:0] w774;
	wire [0:0] w775;
	wire [0:0] w776;
	wire [0:0] w777;
	wire [0:0] w778;
	wire [5:0] w779;
	wire [6:0] w780;
	wire [0:0] w781;
	wire [0:0] w782;
	wire [0:0] w783;
	wire [0:0] w785;
	wire [0:0] w786;
	wire [0:0] w787;
	wire [0:0] w788;
	wire [0:0] w789;
	wire [0:0] w790;
	wire [6:0] w791;
	wire [7:0] w794;
	wire [7:0] w795;
	wire [7:0] w796;
	wire [7:0] w799;
	wire [0:0] w800;
	wire [0:0] w801;
	wire [0:0] w802;
	wire [0:0] w803;
	wire [0:0] w804;
	wire [0:0] w805;
	wire [0:0] w806;
	wire [0:0] w807;
	wire [0:0] w808;
	wire [0:0] w809;
	wire [0:0] w810;
	wire [0:0] w811;
	wire [0:0] w812;
	wire [31:0] w814;
	wire [31:0] w816;
	wire [31:0] w817;
	wire [0:0] w818;
	wire [31:0] w819;
	wire [0:0] w820;
	wire [0:0] w821;
	wire [0:0] w822;
	wire [0:0] w823;
	wire [10:0] w824;
	wire [11:0] w825;
	wire [0:0] w826;
	wire [10:0] w827;
	wire [11:0] w828;
	wire [0:0] w829;
	wire [10:0] w830;
	wire [11:0] w831;
	wire [0:0] w832;
	wire [10:0] w833;
	wire [11:0] w834;
	wire [0:0] w835;
	wire [1:0] w836;
	wire [2:0] w837;
	wire [3:0] w838;
	wire [0:0] w839;
	wire [0:0] w840;
	wire [0:0] w841;
	wire [0:0] w842;
	wire [9:0] w843;
	wire [11:0] w844;
	wire [0:0] w845;
	wire [9:0] w846;
	wire [11:0] w847;
	wire [0:0] w848;
	wire [9:0] w849;
	wire [11:0] w850;
	wire [0:0] w851;
	wire [7:0] w852;
	wire [11:0] w853;
	wire [0:0] w854;
	wire [9:0] w855;
	wire [11:0] w856;
	wire [0:0] w857;
	wire [11:0] w858;
	wire [0:0] w859;
	wire [1:0] w860;
	wire [2:0] w861;
	wire [3:0] w862;
	wire [4:0] w863;
	wire [5:0] w864;
	wire [6:0] w865;
	wire [7:0] w866;
	wire [8:0] w867;
	wire [9:0] w868;
	wire [10:0] w869;
	wire [11:0] w870;
	wire [12:0] w871;
	wire [13:0] w873;
	wire [14:0] w875;
	wire [15:0] w876;
	wire [16:0] w878;
	wire [17:0] w880;
	wire [18:0] w882;
	wire [0:0] w883;
	wire [0:0] w884;
	wire [0:0] w886;
	wire [0:0] w887;
	wire [0:0] w888;
	wire [0:0] w889;
	wire [0:0] w890;
	wire [0:0] w891;
	wire [31:0] w892;
	wire [31:0] w893;
	wire [31:0] w894;
	wire [31:0] w895;
	wire [0:0] w897;
	wire [0:0] w899;
	wire [0:0] w901;
	wire [0:0] w902;
	wire [0:0] w903;
	wire [0:0] w904;
	wire [0:0] w905;
	wire [0:0] w906;
	wire [0:0] w907;
	wire [0:0] w908;
	wire [0:0] w909;
	wire [0:0] w910;
	wire [0:0] w911;
	wire [0:0] w912;
	wire [0:0] w913;
	wire [0:0] w914;
	wire [11:0] w915;
	wire [11:0] w916;
	wire [1:0] w918;
	wire [2:0] w919;
	wire [3:0] w920;
	wire [4:0] w921;
	wire [5:0] w922;
	wire [6:0] w923;
	wire [7:0] w924;
	wire [8:0] w925;
	wire [0:0] w926;
	wire [31:0] w927;
	wire [1:0] w928;
	wire [2:0] w929;
	wire [3:0] w930;
	wire [4:0] w931;
	wire [5:0] w932;
	wire [6:0] w933;
	wire [7:0] w934;
	wire [8:0] w935;
	wire [9:0] w936;
	wire [10:0] w937;
	wire [11:0] w938;
	wire [12:0] w939;
	wire [13:0] w940;
	wire [14:0] w941;
	wire [15:0] w942;
	wire [0:0] w943;
	wire [31:0] w944;
	wire [0:0] w945;
	wire [0:0] w946;
	wire [0:0] w947;
	wire [0:0] w948;
	wire [0:0] w949;
	wire [0:0] w950;
	wire [0:0] w951;
	wire [0:0] w952;
	wire [0:0] w953;
	wire [0:0] w954;
	wire [0:0] w955;
	wire [0:0] w956;
	wire [0:0] w957;
	wire [0:0] w958;
	wire [0:0] w961;
	wire [1:0] w962;
	wire [0:0] w963;
	wire [0:0] w964;
	wire [0:0] w965;
	wire [0:0] w966;
	wire [0:0] w968;
	wire [0:0] w969;
	wire [0:0] w970;
	wire [1:0] w971;
	wire [0:0] w972;
	wire [0:0] w973;
	wire [1:0] w974;
	wire [0:0] w975;
	wire [0:0] w976;
	wire [0:0] w977;
	wire [0:0] w978;
	wire [0:0] w979;
	wire [0:0] w980;
	wire [0:0] w981;
	wire [0:0] w982;
	wire [0:0] w983;
	wire [31:0] w985;
	wire [0:0] w986;
	wire [3:0] w987;
	wire [0:0] w988;
	wire [31:0] w989;
	wire [1:0] w990;
	wire [0:0] w991;
	wire [31:0] w992;
	wire [0:0] w993;
	wire [0:0] w994;
	wire [0:0] w995;
	wire [0:0] w996;
	wire [0:0] w997;
	wire [2:0] w998;
	wire [31:0] w999;
	wire [0:0] w1000;
	wire [0:0] w1001;
	wire [2:0] w1002;
	wire [31:0] w1003;
	wire [63:0] w1005;
	wire [63:0] w1006;
	wire [63:0] w1010;
	wire [31:0] w1013;
	wire [31:0] w1014;
	wire [31:0] w1015;
	wire [31:0] w1016;
	wire [31:0] w1017;
	wire [9:0] w1018;
	wire [11:0] w1019;
	wire [0:0] w1020;
	wire [31:0] w1021;
	wire [31:0] w1022;
	wire [31:0] w1023;
	wire [31:0] w1024;
	wire [6:0] w1025;
	wire [0:0] w1026;
	wire [31:0] w1027;
	wire [31:0] w1028;
	wire [31:0] w1029;
	wire [31:0] w1030;
	wire [31:0] w1031;
	wire [31:0] w1032;
	wire [11:0] w1033;
	wire [31:0] w1034;
	wire [0:0] w1035;
	wire [31:0] w1036;
	wire [31:0] w1037;
	wire [11:0] w1038;
	wire [31:0] w1039;
	wire [0:0] w1040;
	wire [31:0] w1041;
	wire [63:0] w1042;
	wire [31:0] w1045;
	wire [11:0] w1046;
	wire [31:0] w1047;
	wire [0:0] w1048;
	wire [31:0] w1049;
	wire [31:0] w1050;
	wire [11:0] w1051;
	wire [31:0] w1052;
	wire [0:0] w1053;
	wire [31:0] w1054;
	wire [31:0] w1055;
	wire [11:0] w1056;
	wire [31:0] w1057;
	wire [0:0] w1058;
	wire [31:0] w1059;
	wire [31:0] w1060;
	wire [11:0] w1061;
	wire [31:0] w1062;
	wire [0:0] w1063;
	wire [31:0] w1064;
	wire [31:0] w1065;
	wire [31:0] w1067;
	wire [31:0] w1068;
	wire [0:0] w1071;
	wire [0:0] w1072;
	wire [0:0] w1073;
	wire [31:0] w1074;
	wire [0:0] w1075;
	wire [31:0] w1076;
	wire [31:0] w1077;
	wire [0:0] w1078;
	wire [0:0] w1079;
	wire [11:0] w1080;
	wire [31:0] w1081;
	wire [31:0] w1082;
	wire [31:0] w1083;
	wire [31:0] w1084;
	wire [1:0] w1085;
	wire [0:0] w1086;
	wire [31:0] w1087;
	wire [31:0] w1088;
	wire [31:0] w1089;
	wire [31:0] w1090;
	wire [0:0] w1091;
	wire [0:0] w1092;
	wire [0:0] w1093;
	wire [0:0] w1094;
	wire [0:0] w1095;
	wire [0:0] w1096;
	wire [0:0] w1097;
	wire [0:0] w1098;
	wire [0:0] w1099;
	wire [0:0] w1100;
	wire [0:0] w1101;
	wire [0:0] w1102;
	wire [0:0] w1103;
	wire [0:0] w1104;
	wire [0:0] w1105;
	wire [0:0] w1106;
	wire [31:0] w1107;
	wire [0:0] w1108;
	wire [4:0] w1109;
	wire [4:0] w1110;
	wire [4:0] w1111;
	wire [4:0] w1112;
	wire [0:0] w1113;
	wire [31:0] w1114;
	wire [0:0] w1115;
	wire [31:0] w1116;
	wire [31:0] w1117;
	wire [31:0] w1118;
	wire [4:0] w1119;
	wire [0:0] w1120;
	wire [31:0] w1121;
	wire [4:0] w1122;
	wire [31:0] w1123;
	wire [4:0] w1124;
	wire [0:0] w1125;
	wire [0:0] w1126;
	wire [0:0] w1128;
	wire [0:0] w1130;
	wire [1:0] w1131;
	wire [0:0] w1132;
	wire [1:0] w1133;
	wire [0:0] w1135;
	wire [0:0] w1136;
	wire [1:0] w1137;
	wire [0:0] w1138;
	wire [1:0] w1139;
	wire [1:0] w1140;
	wire [0:0] w1141;
	wire [1:0] w1142;
	wire [0:0] w1143;
	wire [1:0] w1144;
	wire [0:0] w1145;
	wire [0:0] w1146;
	wire [1:0] w1147;
	wire [1:0] w1148;
	wire [4:0] w1149;
	wire [0:0] w1150;
	wire [2:0] w1151;
	wire [2:0] w1152;
	wire [2:0] w1153;
	wire [2:0] w1154;
	wire [0:0] w1155;
	wire [0:0] w1156;
	wire [0:0] w1157;
	wire [33:0] w1161;
	wire [33:0] w1162;
	wire [0:0] w1163;
	wire [33:0] w1164;
	wire [33:0] w1165;
	wire [30:0] w1167;
	wire [31:0] w1168;
	wire [31:0] w1169;
	wire [31:0] w1170;
	wire [31:0] w1171;
	wire [0:0] w1172;
	wire [31:0] w1173;
	wire [31:0] w1174;
	wire [15:0] w1175;
	wire [16:0] w1176;
	wire [16:0] w1177;
	wire [30:0] w1178;
	wire [31:0] w1179;
	wire [31:0] w1180;
	wire [31:0] w1181;
	wire [31:0] w1182;
	wire [0:0] w1183;
	wire [31:0] w1184;
	wire [1:0] w1185;
	wire [0:0] w1186;
	wire [31:0] w1187;
	wire [15:0] w1188;
	wire [16:0] w1189;
	wire [16:0] w1190;
	wire [16:0] w1192;
	wire [16:0] w1193;
	wire [16:0] w1194;
	wire [16:0] w1195;
	wire [0:0] w1196;
	wire [0:0] w1197;
	wire [0:0] w1198;
	wire [0:0] w1199;
	wire [0:0] w1200;
	wire [0:0] w1202;
	wire [1:0] w1204;
	wire [0:0] w1205;
	wire [1:0] w1206;
	wire [4:0] w1208;
	wire [0:0] w1209;
	wire [0:0] w1210;
	wire [1:0] w1211;
	wire [0:0] w1212;
	wire [1:0] w1213;
	wire [1:0] w1214;
	wire [0:0] w1215;
	wire [1:0] w1216;
	wire [0:0] w1217;
	wire [1:0] w1218;
	wire [0:0] w1219;
	wire [0:0] w1220;
	wire [1:0] w1221;
	wire [1:0] w1222;
	wire [4:0] w1223;
	wire [0:0] w1224;
	wire [2:0] w1225;
	wire [2:0] w1226;
	wire [2:0] w1227;
	wire [2:0] w1228;
	wire [0:0] w1229;
	wire [0:0] w1230;
	wire [0:0] w1231;
	wire [35:0] w1235;
	wire [35:0] w1236;
	wire [0:0] w1237;
	wire [35:0] w1238;
	wire [35:0] w1239;
	wire [15:0] w1240;
	wire [16:0] w1241;
	wire [15:0] w1242;
	wire [16:0] w1243;
	wire [16:0] w1244;
	wire [17:0] w1245;
	wire [17:0] w1246;
	wire [15:0] w1247;
	wire [16:0] w1248;
	wire [15:0] w1249;
	wire [16:0] w1250;
	wire [16:0] w1251;
	wire [17:0] w1252;
	wire [17:0] w1253;
	wire [17:0] w1255;
	wire [17:0] w1256;
	wire [17:0] w1257;
	wire [17:0] w1258;
	wire [0:0] w1259;
	wire [0:0] w1260;
	wire [0:0] w1261;
	wire [0:0] w1262;
	wire [0:0] w1263;
	wire [0:0] w1265;
	wire [1:0] w1267;
	wire [0:0] w1268;
	wire [1:0] w1269;
	wire [0:0] w1271;
	wire [0:0] w1272;
	wire [1:0] w1273;
	wire [0:0] w1274;
	wire [1:0] w1275;
	wire [1:0] w1276;
	wire [0:0] w1277;
	wire [1:0] w1278;
	wire [0:0] w1279;
	wire [1:0] w1280;
	wire [0:0] w1281;
	wire [0:0] w1282;
	wire [1:0] w1283;
	wire [1:0] w1284;
	wire [4:0] w1285;
	wire [0:0] w1286;
	wire [2:0] w1287;
	wire [2:0] w1288;
	wire [2:0] w1289;
	wire [2:0] w1290;
	wire [0:0] w1291;
	wire [0:0] w1292;
	wire [0:0] w1293;
	wire [33:0] w1295;
	wire [0:0] w1296;
	wire [33:0] w1297;
	wire [33:0] w1298;
	wire [15:0] w1299;
	wire [16:0] w1300;
	wire [16:0] w1301;
	wire [15:0] w1302;
	wire [16:0] w1303;
	wire [16:0] w1304;
	wire [16:0] w1306;
	wire [16:0] w1307;
	wire [16:0] w1308;
	wire [16:0] w1309;
	wire [0:0] w1310;
	wire [0:0] w1311;
	wire [0:0] w1312;
	wire [0:0] w1313;
	wire [0:0] w1314;
	wire [0:0] w1315;
	wire [0:0] w1316;
	wire [17:0] w1317;
	wire [17:0] w1318;
	wire [35:0] w1319;
	wire [35:0] w1320;
	wire [35:0] w1321;
	wire [35:0] w1322;
	wire [35:0] w1323;
	wire [35:0] w1324;
	wire [31:0] w1325;
	wire [63:0] w1326;
	wire [35:0] w1327;
	wire [35:0] w1328;
	wire [51:0] w1330;
	wire [0:0] w1331;
	wire [52:0] w1333;
	wire [0:0] w1334;
	wire [53:0] w1336;
	wire [0:0] w1337;
	wire [54:0] w1339;
	wire [0:0] w1340;
	wire [55:0] w1342;
	wire [0:0] w1343;
	wire [56:0] w1345;
	wire [0:0] w1346;
	wire [57:0] w1348;
	wire [0:0] w1349;
	wire [58:0] w1351;
	wire [0:0] w1352;
	wire [59:0] w1354;
	wire [0:0] w1355;
	wire [60:0] w1357;
	wire [0:0] w1358;
	wire [61:0] w1360;
	wire [0:0] w1361;
	wire [62:0] w1363;
	wire [0:0] w1364;
	wire [63:0] w1365;
	wire [63:0] w1366;
	wire [0:0] w1367;
	wire [34:0] w1368;
	wire [0:0] w1369;
	wire [35:0] w1370;
	wire [0:0] w1371;
	wire [36:0] w1372;
	wire [0:0] w1373;
	wire [37:0] w1375;
	wire [0:0] w1376;
	wire [38:0] w1378;
	wire [0:0] w1379;
	wire [39:0] w1381;
	wire [0:0] w1382;
	wire [40:0] w1384;
	wire [0:0] w1385;
	wire [41:0] w1387;
	wire [0:0] w1388;
	wire [42:0] w1390;
	wire [0:0] w1391;
	wire [43:0] w1393;
	wire [0:0] w1394;
	wire [44:0] w1396;
	wire [0:0] w1397;
	wire [45:0] w1399;
	wire [0:0] w1400;
	wire [46:0] w1402;
	wire [0:0] w1403;
	wire [47:0] w1405;
	wire [0:0] w1406;
	wire [48:0] w1408;
	wire [0:0] w1409;
	wire [49:0] w1411;
	wire [0:0] w1412;
	wire [50:0] w1414;
	wire [0:0] w1415;
	wire [51:0] w1416;
	wire [0:0] w1417;
	wire [52:0] w1418;
	wire [0:0] w1419;
	wire [53:0] w1420;
	wire [0:0] w1421;
	wire [54:0] w1422;
	wire [0:0] w1423;
	wire [55:0] w1424;
	wire [0:0] w1425;
	wire [56:0] w1426;
	wire [0:0] w1427;
	wire [57:0] w1428;
	wire [0:0] w1429;
	wire [58:0] w1430;
	wire [0:0] w1431;
	wire [59:0] w1432;
	wire [0:0] w1433;
	wire [60:0] w1434;
	wire [0:0] w1435;
	wire [61:0] w1436;
	wire [0:0] w1437;
	wire [62:0] w1438;
	wire [0:0] w1439;
	wire [63:0] w1440;
	wire [63:0] w1441;
	wire [63:0] w1442;
	wire [63:0] w1443;
	wire [63:0] w1444;
	wire [63:0] w1445;
	wire [2:0] w1446;
	wire [2:0] w1447;
	wire [2:0] w1448;
	wire [0:0] w1449;
	wire [0:0] w1450;
	wire [0:0] w1451;
	wire [0:0] w1452;
	wire [0:0] w1453;
	wire [0:0] w1454;
	wire [15:0] w1455;
	wire [15:0] w1456;
	wire [15:0] w1457;
	wire [15:0] w1458;
	wire [33:0] w1459;
	wire [35:0] w1460;
	wire [35:0] w1461;
	wire [33:0] w1462;
	wire [0:0] w1463;
	wire [11:0] w1464;
	wire [0:0] w1465;
	wire [31:0] w1466;
	wire [0:0] w1468;
	wire [31:0] w1469;
	wire [31:0] w1470;
	wire [0:0] w1471;
	wire [0:0] w1472;
	wire [0:0] w1473;
	wire [0:0] w1474;
	wire [31:0] w1476;
	wire [31:0] w1477;
	wire [31:0] w1478;
	wire [1:0] w1479;
	wire [2:0] w1480;
	wire [0:0] w1481;
	wire [31:0] w1482;
	wire [31:0] w1483;
	wire [31:0] w1484;
	wire [16:0] w1485;
	wire [31:0] w1486;
	wire [16:0] w1487;
	wire [0:0] w1488;
	wire [0:0] w1489;
	wire [0:0] w1494;
	wire [31:0] w1495;
	wire [31:0] w1498;
	wire [0:0] w1499;
	wire [31:0] w1500;
	wire [31:0] w1503;
	wire [31:0] w1506;
	wire [31:0] w1507;
	wire [0:0] w1508;
	wire [31:0] w1509;
	wire [31:0] w1512;
	wire [31:0] w1515;
	wire [31:0] w1516;
	wire [31:0] w1519;
	wire [31:0] w1522;
	wire [31:0] w1523;
	wire [31:0] w1524;
	wire [0:0] w1525;
	wire [31:0] w1526;
	wire [31:0] w1529;
	wire [31:0] w1532;
	wire [31:0] w1533;
	wire [31:0] w1536;
	wire [31:0] w1539;
	wire [31:0] w1540;
	wire [31:0] w1541;
	wire [31:0] w1544;
	wire [31:0] w1547;
	wire [31:0] w1548;
	wire [31:0] w1551;
	wire [31:0] w1554;
	wire [31:0] w1555;
	wire [31:0] w1556;
	wire [31:0] w1557;
	wire [0:0] w1558;
	wire [31:0] w1559;
	wire [31:0] w1562;
	wire [31:0] w1565;
	wire [31:0] w1566;
	wire [31:0] w1569;
	wire [31:0] w1572;
	wire [31:0] w1573;
	wire [31:0] w1574;
	wire [31:0] w1577;
	wire [31:0] w1580;
	wire [31:0] w1581;
	wire [31:0] w1584;
	wire [31:0] w1587;
	wire [31:0] w1588;
	wire [31:0] w1589;
	wire [31:0] w1590;
	wire [31:0] w1593;
	wire [31:0] w1596;
	wire [31:0] w1597;
	wire [31:0] w1600;
	wire [31:0] w1603;
	wire [31:0] w1604;
	wire [31:0] w1605;
	wire [31:0] w1608;
	wire [31:0] w1611;
	wire [31:0] w1612;
	wire [31:0] w1615;
	wire [31:0] w1618;
	wire [31:0] w1619;
	wire [31:0] w1620;
	wire [31:0] w1621;
	wire [31:0] w1622;
	wire [0:0] w1623;
	wire [31:0] w1624;
	wire [31:0] w1627;
	wire [31:0] w1630;
	wire [31:0] w1631;
	wire [31:0] w1634;
	wire [31:0] w1637;
	wire [31:0] w1638;
	wire [31:0] w1639;
	wire [31:0] w1642;
	wire [31:0] w1645;
	wire [31:0] w1646;
	wire [31:0] w1649;
	wire [31:0] w1652;
	wire [31:0] w1653;
	wire [31:0] w1654;
	wire [31:0] w1655;
	wire [31:0] w1658;
	wire [31:0] w1661;
	wire [31:0] w1662;
	wire [31:0] w1665;
	wire [31:0] w1668;
	wire [31:0] w1669;
	wire [31:0] w1670;
	wire [31:0] w1673;
	wire [31:0] w1676;
	wire [31:0] w1677;
	wire [31:0] w1680;
	wire [31:0] w1683;
	wire [31:0] w1684;
	wire [31:0] w1685;
	wire [31:0] w1686;
	wire [31:0] w1687;
	wire [31:0] w1690;
	wire [31:0] w1693;
	wire [31:0] w1694;
	wire [31:0] w1697;
	wire [31:0] w1700;
	wire [31:0] w1701;
	wire [31:0] w1702;
	wire [31:0] w1705;
	wire [31:0] w1708;
	wire [31:0] w1709;
	wire [31:0] w1712;
	wire [31:0] w1715;
	wire [31:0] w1716;
	wire [31:0] w1717;
	wire [31:0] w1718;
	wire [31:0] w1721;
	wire [31:0] w1724;
	wire [31:0] w1725;
	wire [31:0] w1728;
	wire [31:0] w1731;
	wire [31:0] w1732;
	wire [31:0] w1733;
	wire [31:0] w1736;
	wire [31:0] w1739;
	wire [31:0] w1740;
	wire [31:0] w1743;
	wire [31:0] w1746;
	wire [31:0] w1747;
	wire [31:0] w1748;
	wire [31:0] w1749;
	wire [31:0] w1750;
	wire [31:0] w1751;
	wire [0:0] w1752;
	wire [31:0] w1753;
	wire [31:0] w1756;
	wire [31:0] w1759;
	wire [31:0] w1760;
	wire [31:0] w1763;
	wire [31:0] w1766;
	wire [31:0] w1767;
	wire [31:0] w1768;
	wire [31:0] w1771;
	wire [31:0] w1774;
	wire [31:0] w1775;
	wire [31:0] w1778;
	wire [31:0] w1781;
	wire [31:0] w1782;
	wire [31:0] w1783;
	wire [31:0] w1784;
	wire [31:0] w1787;
	wire [31:0] w1790;
	wire [31:0] w1791;
	wire [31:0] w1794;
	wire [31:0] w1797;
	wire [31:0] w1798;
	wire [31:0] w1799;
	wire [31:0] w1802;
	wire [31:0] w1805;
	wire [31:0] w1806;
	wire [31:0] w1809;
	wire [31:0] w1812;
	wire [31:0] w1813;
	wire [31:0] w1814;
	wire [31:0] w1815;
	wire [31:0] w1816;
	wire [31:0] w1819;
	wire [31:0] w1822;
	wire [31:0] w1823;
	wire [31:0] w1826;
	wire [31:0] w1829;
	wire [31:0] w1830;
	wire [31:0] w1831;
	wire [31:0] w1834;
	wire [31:0] w1837;
	wire [31:0] w1838;
	wire [31:0] w1841;
	wire [31:0] w1844;
	wire [31:0] w1845;
	wire [31:0] w1846;
	wire [31:0] w1847;
	wire [31:0] w1850;
	wire [31:0] w1853;
	wire [31:0] w1854;
	wire [31:0] w1857;
	wire [31:0] w1860;
	wire [31:0] w1861;
	wire [31:0] w1862;
	wire [31:0] w1865;
	wire [31:0] w1868;
	wire [31:0] w1869;
	wire [31:0] w1872;
	wire [31:0] w1875;
	wire [31:0] w1876;
	wire [31:0] w1877;
	wire [31:0] w1878;
	wire [31:0] w1879;
	wire [31:0] w1880;
	wire [31:0] w1883;
	wire [31:0] w1886;
	wire [31:0] w1887;
	wire [31:0] w1890;
	wire [31:0] w1893;
	wire [31:0] w1894;
	wire [31:0] w1895;
	wire [31:0] w1898;
	wire [31:0] w1901;
	wire [31:0] w1902;
	wire [31:0] w1905;
	wire [31:0] w1908;
	wire [31:0] w1909;
	wire [31:0] w1910;
	wire [31:0] w1911;
	wire [31:0] w1914;
	wire [31:0] w1917;
	wire [31:0] w1918;
	wire [31:0] w1921;
	wire [31:0] w1924;
	wire [31:0] w1925;
	wire [31:0] w1926;
	wire [31:0] w1929;
	wire [31:0] w1932;
	wire [31:0] w1933;
	wire [31:0] w1936;
	wire [31:0] w1939;
	wire [31:0] w1940;
	wire [31:0] w1941;
	wire [31:0] w1942;
	wire [31:0] w1943;
	wire [31:0] w1946;
	wire [31:0] w1949;
	wire [31:0] w1950;
	wire [31:0] w1953;
	wire [31:0] w1956;
	wire [31:0] w1957;
	wire [31:0] w1958;
	wire [31:0] w1961;
	wire [31:0] w1964;
	wire [31:0] w1965;
	wire [31:0] w1968;
	wire [31:0] w1971;
	wire [31:0] w1972;
	wire [31:0] w1973;
	wire [31:0] w1974;
	wire [31:0] w1977;
	wire [31:0] w1980;
	wire [31:0] w1981;
	wire [31:0] w1984;
	wire [31:0] w1987;
	wire [31:0] w1988;
	wire [31:0] w1989;
	wire [31:0] w1992;
	wire [31:0] w1995;
	wire [31:0] w1996;
	wire [31:0] w1999;
	wire [31:0] w2002;
	wire [31:0] w2003;
	wire [31:0] w2004;
	wire [31:0] w2005;
	wire [31:0] w2006;
	wire [31:0] w2007;
	wire [31:0] w2008;
	wire [31:0] w2009;
	wire [31:0] w2010;
	wire [30:0] w2011;
	wire [31:0] w2012;
	wire [31:0] w2013;
	wire [4:0] w2014;
	wire [4:0] w2015;
	wire [0:0] w2016;
	wire [4:0] w2017;
	wire [4:0] w2018;
	wire [4:0] w2019;
	wire [4:0] w2020;
	wire [4:0] w2021;
	wire [31:0] w2022;
	wire [3:0] w2023;
	wire [4:0] w2024;
	wire [0:0] w2025;
	wire [0:0] w2026;
	wire [4:0] w2027;
	wire [3:0] w2028;
	wire [4:0] w2029;
	wire [0:0] w2030;
	wire [0:0] w2031;
	wire [4:0] w2032;
	wire [1:0] w2033;
	wire [14:0] w2034;
	wire [19:0] w2036;
	wire [24:0] w2038;
	wire [4:0] w2039;
	wire [29:0] w2041;
	wire [31:0] w2042;
	wire [6:0] w2043;
	wire [6:0] w2044;
	wire [0:0] w2045;
	wire [2:0] w2046;
	wire [2:0] w2047;
	wire [0:0] w2048;
	wire [0:0] w2049;
	wire [31:0] w2050;
	wire [3:0] w2051;
	wire [4:0] w2052;
	wire [0:0] w2053;
	wire [0:0] w2054;
	wire [4:0] w2055;
	wire [6:0] w2056;
	wire [11:0] w2057;
	wire [2:0] w2058;
	wire [14:0] w2059;
	wire [19:0] w2060;
	wire [9:0] w2061;
	wire [29:0] w2062;
	wire [31:0] w2063;
	wire [6:0] w2064;
	wire [0:0] w2065;
	wire [0:0] w2066;
	wire [31:0] w2067;
	wire [6:0] w2068;
	wire [11:0] w2069;
	wire [2:0] w2070;
	wire [14:0] w2071;
	wire [19:0] w2072;
	wire [11:0] w2073;
	wire [31:0] w2074;
	wire [6:0] w2075;
	wire [0:0] w2076;
	wire [31:0] w2077;
	wire [6:0] w2078;
	wire [11:0] w2079;
	wire [2:0] w2080;
	wire [14:0] w2081;
	wire [19:0] w2082;
	wire [24:0] w2083;
	wire [6:0] w2084;
	wire [31:0] w2085;
	wire [6:0] w2086;
	wire [0:0] w2087;
	wire [31:0] w2088;
	wire [31:0] w2089;
	wire [31:0] w2090;
	wire [6:0] w2091;
	wire [6:0] w2092;
	wire [6:0] w2093;
	wire [4:0] w2094;
	wire [11:0] w2095;
	wire [11:0] w2096;
	wire [31:0] w2097;
	wire [6:0] w2098;
	wire [2:0] w2099;
	wire [0:0] w2100;
	wire [0:0] w2101;
	wire [0:0] w2102;
	wire [0:0] w2103;
	wire [0:0] w2104;
	wire [0:0] w2105;
	wire [0:0] w2106;
	wire [0:0] w2107;
	wire [0:0] w2108;
	wire [0:0] w2109;
	wire [0:0] w2110;
	wire [31:0] w2111;
	wire [0:0] w2112;
	wire [31:0] w2113;
	wire [0:0] w2114;
	wire [0:0] w2115;
	wire [0:0] w2116;
	wire [31:0] w2117;
	wire [0:0] w2118;
	wire [0:0] w2119;
	wire [31:0] w2120;
	wire [6:0] w2121;
	wire [11:0] w2122;
	wire [2:0] w2123;
	wire [14:0] w2124;
	wire [19:0] w2125;
	wire [9:0] w2126;
	wire [29:0] w2127;
	wire [29:0] w2128;
	wire [31:0] w2129;
	wire [14:0] w2130;
	wire [19:0] w2131;
	wire [24:0] w2132;
	wire [4:0] w2133;
	wire [29:0] w2134;
	wire [29:0] w2135;
	wire [0:0] w2136;
	wire [0:0] w2137;
	wire [0:0] w2138;
	wire [0:0] w2139;
	wire [9:0] w2140;
	wire [9:0] w2141;
	wire [4:0] w2142;
	wire [4:0] w2143;
	wire [4:0] w2144;
	wire [4:0] w2145;
	wire [4:0] w2146;
	wire [2:0] w2147;
	wire [6:0] w2148;
	wire [11:0] w2149;
	wire [4:0] w2150;
	wire [6:0] w2151;
	wire [6:0] w2152;
	wire [31:0] w2153;
	wire [31:0] w2154;
	wire [4:0] w2155;
	wire [4:0] w2156;
	wire [4:0] w2157;
	wire [4:0] w2158;
	wire [0:0] w2159;
	wire [0:0] w2160;
	wire [31:0] w2161;
	wire [31:0] w2162;
	wire [0:0] w2163;
	wire [0:0] w2164;
	wire [0:0] w2165;
	wire [0:0] w2166;
	wire [2:0] w2167;
	wire [6:0] w2168;
	wire [31:0] w2169;
	wire [11:0] w2170;
	wire [4:0] w2171;
	wire [6:0] w2172;
	wire [6:0] w2173;
	wire [4:0] w2174;
	wire [4:0] w2175;
	wire [4:0] w2176;
	wire [4:0] w2177;
	wire [31:0] w2178;
	wire [0:0] w2179;
	wire [0:0] w2180;
	wire [31:0] w2181;
	wire [0:0] w2182;
	wire [0:0] w2183;
	wire [0:0] w2184;
	wire [0:0] w2185;
	wire [0:0] w2186;
	wire [31:0] w2187;
	wire [0:0] w2192;
	wire [0:0] w2193;
	wire [1:0] w2194;
	wire [0:0] w2195;
	wire [2:0] w2196;
	wire [0:0] w2197;
	wire [3:0] w2198;
	wire [0:0] w2199;
	wire [4:0] w2200;
	wire [0:0] w2201;
	wire [5:0] w2202;
	wire [0:0] w2203;
	wire [6:0] w2204;
	wire [0:0] w2205;
	wire [7:0] w2206;
	wire [0:0] w2207;
	wire [8:0] w2208;
	wire [0:0] w2209;
	wire [9:0] w2210;
	wire [0:0] w2211;
	wire [10:0] w2212;
	wire [0:0] w2213;
	wire [11:0] w2214;
	wire [0:0] w2215;
	wire [12:0] w2216;
	wire [0:0] w2217;
	wire [13:0] w2218;
	wire [0:0] w2219;
	wire [14:0] w2220;
	wire [0:0] w2221;
	wire [15:0] w2222;
	wire [0:0] w2223;
	wire [16:0] w2224;
	wire [0:0] w2225;
	wire [17:0] w2226;
	wire [0:0] w2227;
	wire [18:0] w2228;
	wire [0:0] w2229;
	wire [19:0] w2230;
	wire [0:0] w2231;
	wire [20:0] w2233;
	wire [0:0] w2234;
	wire [21:0] w2236;
	wire [0:0] w2237;
	wire [22:0] w2239;
	wire [0:0] w2240;
	wire [23:0] w2241;
	wire [23:0] w2242;
	wire [23:0] w2243;
	wire [0:0] w2244;
	wire [23:0] w2245;
	wire [7:0] w2246;
	wire [31:0] w2247;
	wire [0:0] w2248;
	wire [31:0] w2249;
	wire [0:0] w2251;
	wire [0:0] w2252;
	wire [1:0] w2253;
	wire [0:0] w2254;
	wire [2:0] w2255;
	wire [0:0] w2256;
	wire [3:0] w2257;
	wire [0:0] w2258;
	wire [4:0] w2259;
	wire [0:0] w2260;
	wire [5:0] w2261;
	wire [0:0] w2262;
	wire [6:0] w2263;
	wire [0:0] w2264;
	wire [7:0] w2265;
	wire [0:0] w2266;
	wire [8:0] w2267;
	wire [0:0] w2268;
	wire [9:0] w2269;
	wire [0:0] w2270;
	wire [10:0] w2271;
	wire [0:0] w2272;
	wire [11:0] w2273;
	wire [0:0] w2274;
	wire [12:0] w2275;
	wire [0:0] w2276;
	wire [13:0] w2277;
	wire [0:0] w2278;
	wire [14:0] w2279;
	wire [0:0] w2280;
	wire [15:0] w2281;
	wire [0:0] w2282;
	wire [16:0] w2283;
	wire [0:0] w2284;
	wire [17:0] w2285;
	wire [0:0] w2286;
	wire [18:0] w2287;
	wire [0:0] w2288;
	wire [19:0] w2289;
	wire [0:0] w2290;
	wire [20:0] w2291;
	wire [0:0] w2292;
	wire [21:0] w2293;
	wire [0:0] w2294;
	wire [22:0] w2295;
	wire [0:0] w2296;
	wire [23:0] w2297;
	wire [23:0] w2298;
	wire [23:0] w2299;
	wire [7:0] w2300;
	wire [31:0] w2301;
	wire [0:0] w2302;
	wire [31:0] w2303;
	wire [0:0] w2305;
	wire [0:0] w2306;
	wire [1:0] w2307;
	wire [0:0] w2308;
	wire [2:0] w2309;
	wire [0:0] w2310;
	wire [3:0] w2311;
	wire [0:0] w2312;
	wire [4:0] w2313;
	wire [0:0] w2314;
	wire [5:0] w2315;
	wire [0:0] w2316;
	wire [6:0] w2317;
	wire [0:0] w2318;
	wire [7:0] w2319;
	wire [0:0] w2320;
	wire [8:0] w2321;
	wire [0:0] w2322;
	wire [9:0] w2323;
	wire [0:0] w2324;
	wire [10:0] w2325;
	wire [0:0] w2326;
	wire [11:0] w2327;
	wire [0:0] w2328;
	wire [12:0] w2329;
	wire [0:0] w2330;
	wire [13:0] w2331;
	wire [0:0] w2332;
	wire [14:0] w2333;
	wire [0:0] w2334;
	wire [15:0] w2335;
	wire [0:0] w2336;
	wire [16:0] w2337;
	wire [0:0] w2338;
	wire [17:0] w2339;
	wire [0:0] w2340;
	wire [18:0] w2341;
	wire [0:0] w2342;
	wire [19:0] w2343;
	wire [0:0] w2344;
	wire [20:0] w2345;
	wire [0:0] w2346;
	wire [21:0] w2347;
	wire [0:0] w2348;
	wire [22:0] w2349;
	wire [0:0] w2350;
	wire [23:0] w2351;
	wire [23:0] w2352;
	wire [23:0] w2353;
	wire [7:0] w2354;
	wire [31:0] w2355;
	wire [1:0] w2356;
	wire [0:0] w2357;
	wire [31:0] w2358;
	wire [0:0] w2360;
	wire [0:0] w2361;
	wire [1:0] w2362;
	wire [0:0] w2363;
	wire [2:0] w2364;
	wire [0:0] w2365;
	wire [3:0] w2366;
	wire [0:0] w2367;
	wire [4:0] w2368;
	wire [0:0] w2369;
	wire [5:0] w2370;
	wire [0:0] w2371;
	wire [6:0] w2372;
	wire [0:0] w2373;
	wire [7:0] w2374;
	wire [0:0] w2375;
	wire [8:0] w2376;
	wire [0:0] w2377;
	wire [9:0] w2378;
	wire [0:0] w2379;
	wire [10:0] w2380;
	wire [0:0] w2381;
	wire [11:0] w2382;
	wire [0:0] w2383;
	wire [12:0] w2384;
	wire [0:0] w2385;
	wire [13:0] w2386;
	wire [0:0] w2387;
	wire [14:0] w2388;
	wire [0:0] w2389;
	wire [15:0] w2390;
	wire [0:0] w2391;
	wire [16:0] w2392;
	wire [0:0] w2393;
	wire [17:0] w2394;
	wire [0:0] w2395;
	wire [18:0] w2396;
	wire [0:0] w2397;
	wire [19:0] w2398;
	wire [0:0] w2399;
	wire [20:0] w2400;
	wire [0:0] w2401;
	wire [21:0] w2402;
	wire [0:0] w2403;
	wire [22:0] w2404;
	wire [0:0] w2405;
	wire [23:0] w2406;
	wire [23:0] w2407;
	wire [23:0] w2408;
	wire [7:0] w2409;
	wire [31:0] w2410;
	wire [31:0] w2411;
	wire [0:0] w2412;
	wire [0:0] w2413;
	wire [31:0] w2414;
	wire [15:0] w2417;
	wire [0:0] w2418;
	wire [0:0] w2419;
	wire [1:0] w2420;
	wire [0:0] w2421;
	wire [2:0] w2422;
	wire [0:0] w2423;
	wire [3:0] w2424;
	wire [0:0] w2425;
	wire [4:0] w2426;
	wire [0:0] w2427;
	wire [5:0] w2428;
	wire [0:0] w2429;
	wire [6:0] w2430;
	wire [0:0] w2431;
	wire [7:0] w2432;
	wire [0:0] w2433;
	wire [8:0] w2434;
	wire [0:0] w2435;
	wire [9:0] w2436;
	wire [0:0] w2437;
	wire [10:0] w2438;
	wire [0:0] w2439;
	wire [11:0] w2440;
	wire [0:0] w2441;
	wire [12:0] w2442;
	wire [0:0] w2443;
	wire [13:0] w2444;
	wire [0:0] w2445;
	wire [14:0] w2446;
	wire [0:0] w2447;
	wire [15:0] w2448;
	wire [15:0] w2449;
	wire [15:0] w2450;
	wire [31:0] w2451;
	wire [0:0] w2452;
	wire [31:0] w2453;
	wire [15:0] w2455;
	wire [0:0] w2456;
	wire [0:0] w2457;
	wire [1:0] w2458;
	wire [0:0] w2459;
	wire [2:0] w2460;
	wire [0:0] w2461;
	wire [3:0] w2462;
	wire [0:0] w2463;
	wire [4:0] w2464;
	wire [0:0] w2465;
	wire [5:0] w2466;
	wire [0:0] w2467;
	wire [6:0] w2468;
	wire [0:0] w2469;
	wire [7:0] w2470;
	wire [0:0] w2471;
	wire [8:0] w2472;
	wire [0:0] w2473;
	wire [9:0] w2474;
	wire [0:0] w2475;
	wire [10:0] w2476;
	wire [0:0] w2477;
	wire [11:0] w2478;
	wire [0:0] w2479;
	wire [12:0] w2480;
	wire [0:0] w2481;
	wire [13:0] w2482;
	wire [0:0] w2483;
	wire [14:0] w2484;
	wire [0:0] w2485;
	wire [15:0] w2486;
	wire [15:0] w2487;
	wire [15:0] w2488;
	wire [31:0] w2489;
	wire [0:0] w2490;
	wire [31:0] w2491;
	wire [31:0] w2492;
	wire [31:0] w2493;
	wire [31:0] w2494;
	wire [31:0] w2495;
	wire [31:0] w2496;
	wire [0:0] w2497;
	wire [1:0] w2498;
	wire [1:0] w2500;
	wire [2:0] w2501;
	wire [0:0] w2502;
	wire [31:0] w2503;
	wire [7:0] w2504;
	wire [7:0] w2505;
	wire [15:0] w2506;
	wire [7:0] w2507;
	wire [23:0] w2508;
	wire [7:0] w2509;
	wire [31:0] w2510;
	wire [31:0] w2511;
	wire [15:0] w2512;
	wire [15:0] w2513;
	wire [31:0] w2514;
	wire [31:0] w2515;
	wire [31:0] w2516;
	wire [31:0] w2517;
	wire [31:0] w2518;
	wire [0:0] w2519;
	wire [3:0] w2521;
	wire [3:0] w2522;
	wire [3:0] w2523;
	wire [3:0] w2524;
	wire [3:0] w2525;
	wire [3:0] w2526;
	wire [3:0] w2527;
	wire [3:0] w2528;
	wire [3:0] w2529;
	wire [3:0] w2530;
	wire [3:0] w2531;
	wire [3:0] w2532;
	wire [3:0] w2533;
	wire [0:0] w2534;
	wire [0:0] w2535;
	wire [2:0] w2536;
	wire [2:0] w2537;
	wire [0:0] w2538;
	wire [0:0] w2539;
	wire [0:0] w2540;
	wire [0:0] w2541;
	wire [0:0] w2542;
	wire [0:0] w2543;
	wire [31:0] w2544;
	wire [31:0] w2545;
	wire [3:0] w2546;
	wire [3:0] w2547;
	wire [2:0] w2548;
	wire [3:0] w2549;
	wire [3:0] w2550;
	wire [3:0] w2551;
	wire [2:0] w2552;
	wire [3:0] w2553;
	wire [3:0] w2554;
	wire [3:0] w2555;
	wire [2:0] w2556;
	wire [3:0] w2557;
	wire [3:0] w2558;
	wire [3:0] w2559;
	wire [3:0] w2560;
	wire [3:0] w2561;
	wire [3:0] w2562;
	wire [3:0] w2563;
	wire [1:0] w2564;
	wire [3:0] w2565;
	wire [3:0] w2566;
	wire [0:0] w2567;
	wire [0:0] w2568;
	wire [0:0] w2569;
	wire [1:0] w2570;
	wire [1:0] w2571;
	wire [3:0] w2572;
	wire [3:0] w2573;
	wire [3:0] w2574;
	wire [3:0] w2575;
	wire [3:0] w2576;
	wire [3:0] w2577;
	wire [3:0] w2578;
	wire [3:0] w2579;
	wire [2:0] w2580;
	wire [3:0] w2581;
	wire [3:0] w2582;
	wire [3:0] w2583;
	wire [3:0] w2584;
	wire [3:0] w2585;
	wire [0:0] w2586;
	wire [31:0] w2587;
	wire [0:0] w2588;
	wire [31:0] w2589;
	wire [0:0] w2590;
	wire [0:0] w2591;
	wire [31:0] w2592;
	wire [31:0] w2593;
	wire [0:0] w2594;
	wire [1:0] w2595;
	wire [31:0] w2599;
	wire [0:0] w2603;
	wire [31:0] w2605;
	wire [0:0] w2608;
	wire [0:0] w2610;
	wire [0:0] w2613;
	wire [0:0] w2614;
	wire [0:0] w2616;
	wire [31:0] w2620;
	wire [31:0] w2621;
	wire [0:0] w2622;
	wire [0:0] w2623;
	wire [31:0] w2625;
	wire [0:0] w2628;
	wire [31:0] w2629;
	wire [31:0] w2630;
	wire [0:0] w2631;
	wire [0:0] w2633;
	wire [0:0] w2634;
	wire [0:0] w2635;
	wire [31:0] w2636;
	wire [0:0] w2637;
	wire [0:0] w2638;
	wire [0:0] w2639;
	wire [0:0] w2640;
	wire [0:0] w2641;
	wire [31:0] w2642;
	wire [31:0] w2643;
	wire [31:0] w2644;
	wire [31:0] w2645;
	wire [0:0] w2646;
	wire [8:0] w2647;
	wire [8:0] w2648;
	wire [12:0] w2649;
	wire [5:0] w2650;
	wire [12:0] w2651;
	wire [0:0] w2652;
	wire [8:0] w2653;
	wire [8:0] w2654;
	wire [10:0] w2655;
	wire [12:0] w2656;
	wire [0:0] w2657;
	wire [8:0] w2658;
	wire [8:0] w2659;
	wire [10:0] w2660;
	wire [12:0] w2661;
	wire [0:0] w2662;
	wire [8:0] w2663;
	wire [8:0] w2664;
	wire [10:0] w2665;
	wire [12:0] w2666;
	wire [0:0] w2667;
	wire [8:0] w2668;
	wire [8:0] w2669;
	wire [10:0] w2670;
	wire [12:0] w2671;
	wire [0:0] w2672;
	wire [8:0] w2673;
	wire [8:0] w2674;
	wire [9:0] w2675;
	wire [12:0] w2676;
	wire [0:0] w2677;
	wire [8:0] w2678;
	wire [8:0] w2679;
	wire [9:0] w2680;
	wire [12:0] w2681;
	wire [0:0] w2682;
	wire [8:0] w2683;
	wire [8:0] w2684;
	wire [8:0] w2685;
	wire [12:0] w2686;
	wire [0:0] w2687;
	wire [8:0] w2688;
	wire [8:0] w2689;
	wire [12:0] w2690;
	wire [0:0] w2691;
	wire [8:0] w2692;
	wire [0:0] w2693;
	wire [0:0] w2694;
	wire [0:0] w2695;
	wire [31:0] w2696;
	wire [31:0] w2697;
	wire [11:0] w2698;
	wire [8:0] w2699;
	wire [31:0] w2703;
	wire [31:0] w2704;
	wire [0:0] w2706;
	wire [0:0] w2707;
	wire [0:0] w2708;
	wire [0:0] w2709;
	wire [0:0] w2710;
	wire [0:0] w2711;
	wire [0:0] w2712;
	wire [0:0] w2713;
	wire [0:0] w2714;
	wire [0:0] w2715;
	wire [0:0] w2716;
	wire [0:0] w2717;
	wire [0:0] w2718;
	wire [0:0] w2719;
	wire [0:0] w2720;
	wire [0:0] w2721;
	wire [0:0] w2722;
	wire [31:0] w2723;
	wire [31:0] w2724;
	wire [31:0] w2725;
	wire [31:0] w2726;
	wire [31:0] w2727;
	wire [31:0] w2728;
	wire [31:0] w2730;
	wire [31:0] w2731;
	wire [0:0] w2732;
	wire [0:0] w2733;
	wire [0:0] w2734;
	wire [0:0] w2735;
	wire [0:0] w2736;
	wire [11:0] w2737;
	wire [0:0] w2738;
	wire [0:0] w2739;
	wire [0:0] w2740;
	wire [0:0] w2741;
	wire [0:0] w2742;
	wire [7:0] w2743;
	wire [11:0] w2744;
	wire [0:0] w2745;
	wire [0:0] w2746;
	wire [0:0] w2747;
	wire [6:0] w2748;
	wire [6:0] w2749;
	wire [0:0] w2750;
	wire [6:0] w2751;
	wire [0:0] w2752;
	wire [0:0] w2753;
	wire [0:0] w2754;
	wire [0:0] w2755;
	wire [0:0] w2756;
	wire [0:0] w2757;
	wire [0:0] w2758;
	wire [0:0] w2759;
	wire [1:0] w2761;
	wire [0:0] w2762;
	wire [0:0] w2763;
	wire [0:0] w2764;
	wire [0:0] w2765;
	wire [11:0] w2766;
	wire [31:0] w2767;
	wire [11:0] w2768;
	wire [0:0] w2769;
	wire [12:0] w2770;
	wire [0:0] w2771;
	wire [13:0] w2772;
	wire [0:0] w2773;
	wire [14:0] w2774;
	wire [0:0] w2775;
	wire [15:0] w2776;
	wire [0:0] w2777;
	wire [16:0] w2778;
	wire [0:0] w2779;
	wire [17:0] w2780;
	wire [0:0] w2781;
	wire [18:0] w2782;
	wire [0:0] w2783;
	wire [19:0] w2784;
	wire [0:0] w2785;
	wire [20:0] w2786;
	wire [0:0] w2787;
	wire [21:0] w2788;
	wire [0:0] w2789;
	wire [22:0] w2790;
	wire [0:0] w2791;
	wire [23:0] w2792;
	wire [0:0] w2793;
	wire [24:0] w2794;
	wire [0:0] w2795;
	wire [25:0] w2797;
	wire [0:0] w2798;
	wire [26:0] w2800;
	wire [0:0] w2801;
	wire [27:0] w2803;
	wire [0:0] w2804;
	wire [28:0] w2806;
	wire [0:0] w2807;
	wire [29:0] w2808;
	wire [0:0] w2809;
	wire [30:0] w2810;
	wire [0:0] w2811;
	wire [31:0] w2812;
	wire [31:0] w2813;
	wire [31:0] w2814;
	wire [19:0] w2815;
	wire [11:0] w2816;
	wire [31:0] w2817;
	wire [31:0] w2818;
	wire [31:0] w2819;
	wire [31:0] w2820;
	wire [31:0] w2821;
	wire [31:0] w2822;
	wire [31:0] w2823;
	wire [4:0] w2824;
	wire [6:0] w2825;
	wire [11:0] w2826;
	wire [0:0] w2827;
	wire [12:0] w2828;
	wire [0:0] w2829;
	wire [13:0] w2830;
	wire [0:0] w2831;
	wire [14:0] w2832;
	wire [0:0] w2833;
	wire [15:0] w2834;
	wire [0:0] w2835;
	wire [16:0] w2836;
	wire [0:0] w2837;
	wire [17:0] w2838;
	wire [0:0] w2839;
	wire [18:0] w2840;
	wire [0:0] w2841;
	wire [19:0] w2842;
	wire [0:0] w2843;
	wire [20:0] w2844;
	wire [0:0] w2845;
	wire [21:0] w2846;
	wire [0:0] w2847;
	wire [22:0] w2848;
	wire [0:0] w2849;
	wire [23:0] w2850;
	wire [0:0] w2851;
	wire [24:0] w2852;
	wire [0:0] w2853;
	wire [25:0] w2854;
	wire [0:0] w2855;
	wire [26:0] w2856;
	wire [0:0] w2857;
	wire [27:0] w2858;
	wire [0:0] w2859;
	wire [28:0] w2860;
	wire [0:0] w2861;
	wire [29:0] w2862;
	wire [0:0] w2863;
	wire [30:0] w2864;
	wire [0:0] w2865;
	wire [31:0] w2866;
	wire [31:0] w2867;
	wire [31:0] w2868;
	wire [31:0] w2869;
	wire [31:0] w2870;
	wire [3:0] w2871;
	wire [4:0] w2872;
	wire [5:0] w2873;
	wire [10:0] w2874;
	wire [0:0] w2875;
	wire [11:0] w2876;
	wire [0:0] w2877;
	wire [12:0] w2878;
	wire [0:0] w2879;
	wire [13:0] w2880;
	wire [0:0] w2881;
	wire [14:0] w2882;
	wire [0:0] w2883;
	wire [15:0] w2884;
	wire [0:0] w2885;
	wire [16:0] w2886;
	wire [0:0] w2887;
	wire [17:0] w2888;
	wire [0:0] w2889;
	wire [18:0] w2890;
	wire [0:0] w2891;
	wire [19:0] w2892;
	wire [0:0] w2893;
	wire [20:0] w2894;
	wire [0:0] w2895;
	wire [21:0] w2896;
	wire [0:0] w2897;
	wire [22:0] w2898;
	wire [0:0] w2899;
	wire [23:0] w2900;
	wire [0:0] w2901;
	wire [24:0] w2902;
	wire [0:0] w2903;
	wire [25:0] w2904;
	wire [0:0] w2905;
	wire [26:0] w2906;
	wire [0:0] w2907;
	wire [27:0] w2908;
	wire [0:0] w2909;
	wire [28:0] w2910;
	wire [0:0] w2911;
	wire [29:0] w2912;
	wire [0:0] w2913;
	wire [30:0] w2914;
	wire [0:0] w2915;
	wire [31:0] w2916;
	wire [31:0] w2917;
	wire [31:0] w2918;
	wire [31:0] w2919;
	wire [31:0] w2920;
	wire [9:0] w2921;
	wire [10:0] w2922;
	wire [0:0] w2923;
	wire [11:0] w2924;
	wire [7:0] w2925;
	wire [19:0] w2926;
	wire [0:0] w2927;
	wire [20:0] w2928;
	wire [0:0] w2929;
	wire [21:0] w2930;
	wire [0:0] w2931;
	wire [22:0] w2932;
	wire [0:0] w2933;
	wire [23:0] w2934;
	wire [0:0] w2935;
	wire [24:0] w2936;
	wire [0:0] w2937;
	wire [25:0] w2938;
	wire [0:0] w2939;
	wire [26:0] w2940;
	wire [0:0] w2941;
	wire [27:0] w2942;
	wire [0:0] w2943;
	wire [28:0] w2944;
	wire [0:0] w2945;
	wire [29:0] w2946;
	wire [0:0] w2947;
	wire [30:0] w2948;
	wire [0:0] w2949;
	wire [31:0] w2950;
	wire [31:0] w2951;
	wire [11:0] w2952;
	wire [19:0] w2953;
	wire [31:0] w2954;
	wire [1:0] w2955;
	wire [0:0] w2956;
	wire [31:0] w2957;
	wire [31:0] w2958;
	wire [31:0] w2959;
	wire [4:0] w2960;
	wire [4:0] w2961;
	wire [4:0] w2962;
	wire [31:0] w2963;
	wire [0:0] w2964;
	wire [31:0] w2965;
	wire [0:0] w2966;
	wire [31:0] w2967;
	wire [0:0] w2968;
	wire [31:0] w2969;
	wire [0:0] w2970;
	wire [31:0] w2972;
	wire [0:0] w2973;
	wire [31:0] w2974;
	wire [0:0] w2975;
	wire [0:0] w2976;
	wire [31:0] w2977;
	wire [0:0] w2978;
	wire [31:0] w2979;
	wire [0:0] w2980;
	wire [0:0] w2981;
	wire [31:0] w2982;
	wire [0:0] w2983;
	wire [31:0] w2984;
	wire [0:0] w2985;
	wire [0:0] w2986;
	wire [31:0] w2987;
	wire [0:0] w2988;
	wire [31:0] w2989;
	wire [0:0] w2990;
	wire [31:0] w2992;
	wire [0:0] w2993;
	wire [31:0] w2994;
	wire [0:0] w2996;
	wire [0:0] w2998;
	wire [31:0] w3002;
	wire [0:0] w3003;
	wire [31:0] w3004;
	wire [0:0] w3005;
	wire [31:0] w3007;
	wire [0:0] w3008;
	wire [31:0] w3009;
	wire [0:0] w3010;
	wire [32:0] w3012;
	wire [31:0] w3013;
	wire [0:0] w3014;
	wire [0:0] w3015;
	wire [0:0] w3016;
	wire [0:0] w3017;
	wire [0:0] w3018;
	wire [0:0] w3019;
	wire [31:0] w3020;
	wire [1:0] w3022;
	wire [0:0] w3023;
	wire [31:0] w3024;
	wire [1:0] w3025;
	wire [0:0] w3026;
	wire [31:0] w3027;
	wire [1:0] w3028;
	wire [0:0] w3029;
	wire [31:0] w3030;
	wire [1:0] w3031;
	wire [2:0] w3032;
	wire [3:0] w3033;
	wire [4:0] w3034;
	wire [5:0] w3035;
	wire [0:0] w3036;
	wire [31:0] w3037;
	wire [31:0] w3039;
	wire [1:0] w3042;
	wire [0:0] w3043;
	wire [31:0] w3044;
	wire [31:0] w3046;
	wire [1:0] w3049;
	wire [0:0] w3050;
	wire [31:0] w3051;
	wire [1:0] w3052;
	wire [0:0] w3053;
	wire [31:0] w3054;
	wire [1:0] w3055;
	wire [0:0] w3056;
	wire [31:0] w3057;
	wire [1:0] w3058;
	wire [0:0] w3059;
	wire [31:0] w3060;
	wire [31:0] w3061;
	wire [31:0] w3062;
	wire [31:0] w3063;
	wire [31:0] w3064;
	wire [31:0] w3065;
	wire [31:0] w3066;
	wire [31:0] w3067;
	wire [31:0] w3068;
	wire [31:0] w3069;
	wire [0:0] w3070;
	wire [0:0] w3071;
	wire [0:0] w3072;
	wire [11:0] w3073;
	wire [0:0] w3074;
	wire [31:0] w3075;
	wire [0:0] w3076;
	wire [0:0] w3077;
	wire [0:0] w3078;
	wire [0:0] w3079;
	wire [31:0] w3080;
	wire [31:0] w3081;
	wire [0:0] w3082;
	wire [31:0] w3083;
	wire [31:0] w3084;
	wire [0:0] w3085;
	wire [4:0] w3086;
	wire [4:0] w3087;
	wire [4:0] w3088;
	wire [4:0] w3089;
	wire [6:0] w3090;
	wire [31:0] w3091;
	wire [6:0] w3092;
	wire [4:0] w3093;
	wire [11:0] w3094;
	wire [11:0] w3095;
	wire [6:0] w3096;
	wire [2:0] w3097;
	wire [0:0] w3098;
	wire [0:0] w3099;
	wire [0:0] w3100;
	wire [0:0] w3101;
	wire [0:0] w3102;
	wire [0:0] w3103;
	wire [0:0] w3104;
	wire [0:0] w3105;
	wire [0:0] w3106;
	wire [0:0] w3107;
	wire [0:0] w3108;
	wire [0:0] w3109;
	wire [0:0] w3110;
	wire [0:0] w3111;
	wire [0:0] w3112;
	wire [0:0] w3113;
	wire [0:0] w3114;
	wire [0:0] w3115;
	wire [0:0] w3116;
	wire [0:0] w3117;
	wire [0:0] w3118;
	wire [0:0] w3119;
	wire [0:0] w3120;
	wire [0:0] w3121;
	wire [0:0] w3122;
	wire [0:0] w3123;
	wire [0:0] w3124;
	wire [0:0] w3125;
	wire [0:0] w3126;
	wire [0:0] w3127;
	wire [0:0] w3128;
	wire [0:0] w3129;
	wire [0:0] w3130;
	wire [0:0] w3131;
	wire [0:0] w3132;
	wire [0:0] w3133;
	wire [0:0] w3134;
	wire [31:0] w3135;
	wire [31:0] w3136;
	wire [0:0] w3137;
	wire [31:0] w3138;
	wire [31:0] w3139;
	wire [31:0] w3140;
	wire [31:0] w3141;
	wire [0:0] w3142;
	wire [31:0] w3143;
	wire [31:0] w3144;
	wire [31:0] w3145;
	wire [31:0] w3146;
	wire [31:0] w3147;
	wire [31:0] w3148;
	wire [31:0] w3149;
	wire [31:0] w3150;
	wire [0:0] w3151;
	wire [31:0] w3152;
	wire [31:0] w3153;
	wire [31:0] w3154;
	wire [31:0] w3155;
	wire [31:0] w3156;
	wire [31:0] w3157;
	wire [31:0] w3158;
	wire [31:0] w3159;
	wire [31:0] w3160;
	wire [31:0] w3161;
	wire [31:0] w3162;
	wire [31:0] w3163;
	wire [31:0] w3164;
	wire [31:0] w3165;
	wire [31:0] w3166;
	wire [31:0] w3167;
	wire [0:0] w3168;
	wire [31:0] w3169;
	wire [0:0] w3170;
	wire [31:0] w3171;
	wire [31:0] w3172;
	wire [1:0] w3175;
	wire [3:0] w3176;
	wire [0:0] w3177;
	wire [3:0] w3178;
	wire [0:0] w3179;
	wire [1:0] w3180;
	wire [0:0] w3181;
	wire [1:0] w3182;
	wire [1:0] w3183;
	wire [0:0] w3184;
	wire [1:0] w3185;
	wire [0:0] w3186;
	wire [0:0] w3187;
	wire [1:0] w3188;
	wire [1:0] w3189;
	wire [3:0] w3190;
	wire [0:0] w3191;
	wire [1:0] w3192;
	wire [1:0] w3193;
	wire [0:0] w3194;
	wire [0:0] w3195;
	wire [1:0] w3196;
	wire [1:0] w3197;
	wire [1:0] w3198;
	wire [1:0] w3199;
	wire [31:0] w3201;
	wire [31:0] w3202;
	wire [3:0] w3204;
	wire [0:0] w3206;
	wire [0:0] w3207;
	wire [0:0] w3208;
	wire [0:0] w3209;
	wire [0:0] w3210;
	wire [1:0] w3211;
	wire [0:0] w3212;
	wire [0:0] w3213;
	wire [0:0] w3214;
	wire [0:0] w3215;
	wire [0:0] w3216;
	wire [31:0] w3218;
	wire [3:0] w3220;
	wire [31:0] w3222;
	wire [31:0] w3223;
	wire [31:0] w3224;
	wire [3:0] w3226;
	wire [0:0] w3227;
	wire [0:0] w3228;
	wire [0:0] w3229;
	wire [0:0] w3230;
	wire [0:0] w3231;
	wire [0:0] w3233;
	wire [0:0] w3234;
	wire [0:0] w3237;
	wire [0:0] w3238;
	wire [0:0] w3239;
	wire [0:0] w3240;
	wire [0:0] w3241;
	wire [4:0] w3242;
	wire [0:0] w3243;
	wire [0:0] w3244;
	wire [0:0] w3245;
	wire [0:0] w3246;
	wire [0:0] w3248;
	wire [0:0] w3249;
	wire [3:0] w3250;
	wire [0:0] w3251;
	wire [0:0] w3252;
	wire [0:0] w3253;
	wire [3:0] w3254;
	wire [0:0] w3255;
	wire [0:0] w3256;
	wire [0:0] w3257;
	wire [0:0] w3258;
	wire [0:0] w3259;
	wire [0:0] w3261;
	wire [1:0] w3262;
	wire [0:0] w3263;
	wire [0:0] w3264;
	wire [0:0] w3265;
	wire [1:0] w3266;
	wire [0:0] w3268;
	wire [0:0] w3270;
	wire [0:0] w3271;
	wire [0:0] w3272;
	wire [0:0] w3273;
	wire [0:0] w3274;
	wire [0:0] w3275;
	wire [0:0] w3276;
	wire [0:0] w3277;
	wire [0:0] w3278;
	wire [31:0] w3280;
	wire [15:0] w3282;
	wire [15:0] w3283;
	wire [15:0] w3284;
	wire [15:0] w3286;
	wire [15:0] w3287;
	wire [15:0] w3288;
	wire [31:0] w3292;
	wire [31:0] w3293;
	wire [4:0] w3296;
	wire [4:0] w3297;
	wire [0:0] w3298;
	wire [0:0] w3299;
	wire [0:0] w3300;
	wire [0:0] w3301;
	wire [0:0] w3302;
	wire [0:0] w3303;
	wire [0:0] w3304;
	wire [0:0] w3305;
	wire [0:0] w3306;
	wire [0:0] w3307;
	wire [0:0] w3308;
	wire [0:0] w3309;
	wire [0:0] w3310;
	wire [0:0] w3311;
	wire [0:0] w3312;
	wire [0:0] w3313;
	wire [0:0] w3314;
	wire [31:0] w3315;
	wire [0:0] w3317;
	wire [0:0] w3318;
	wire [0:0] w3319;
	wire [0:0] w3320;
	wire [31:0] w3321;
	wire [0:0] w3323;
	wire [0:0] w3324;
	wire [0:0] w3325;
	wire [0:0] w3326;
	wire [31:0] w3327;
	wire [0:0] w3329;
	wire [0:0] w3330;
	wire [0:0] w3331;
	wire [31:0] w3332;
	wire [0:0] w3334;
	wire [0:0] w3335;
	wire [0:0] w3336;
	wire [0:0] w3337;
	wire [31:0] w3338;
	wire [0:0] w3340;
	wire [0:0] w3341;
	wire [31:0] w3342;
	wire [0:0] w3344;
	wire [0:0] w3345;
	wire [31:0] w3346;
	wire [0:0] w3348;
	wire [0:0] w3349;
	wire [31:0] w3350;
	wire [0:0] w3352;
	wire [0:0] w3353;
	wire [0:0] w3354;
	wire [0:0] w3355;
	wire [0:0] w3356;
	wire [31:0] w3357;
	wire [0:0] w3359;
	wire [0:0] w3360;
	wire [31:0] w3361;
	wire [0:0] w3363;
	wire [0:0] w3364;
	wire [31:0] w3365;
	wire [0:0] w3367;
	wire [0:0] w3368;
	wire [31:0] w3369;
	wire [0:0] w3371;
	wire [0:0] w3372;
	wire [0:0] w3373;
	wire [31:0] w3374;
	wire [0:0] w3376;
	wire [0:0] w3377;
	wire [31:0] w3378;
	wire [0:0] w3380;
	wire [0:0] w3381;
	wire [31:0] w3382;
	wire [0:0] w3384;
	wire [0:0] w3385;
	wire [31:0] w3386;
	wire [0:0] w3388;
	wire [0:0] w3389;
	wire [0:0] w3390;
	wire [0:0] w3391;
	wire [0:0] w3392;
	wire [31:0] w3393;
	wire [0:0] w3395;
	wire [0:0] w3396;
	wire [31:0] w3397;
	wire [0:0] w3399;
	wire [0:0] w3400;
	wire [31:0] w3401;
	wire [0:0] w3403;
	wire [0:0] w3404;
	wire [31:0] w3405;
	wire [0:0] w3407;
	wire [0:0] w3408;
	wire [0:0] w3409;
	wire [31:0] w3410;
	wire [0:0] w3412;
	wire [0:0] w3413;
	wire [31:0] w3414;
	wire [0:0] w3416;
	wire [0:0] w3417;
	wire [31:0] w3418;
	wire [0:0] w3420;
	wire [0:0] w3421;
	wire [31:0] w3422;
	wire [0:0] w3424;
	wire [0:0] w3425;
	wire [0:0] w3426;
	wire [0:0] w3427;
	wire [31:0] w3428;
	wire [0:0] w3430;
	wire [0:0] w3431;
	wire [31:0] w3432;
	wire [0:0] w3434;
	wire [0:0] w3435;
	wire [31:0] w3436;
	wire [0:0] w3438;
	wire [0:0] w3439;
	wire [31:0] w3440;
	wire [0:0] w3442;
	wire [0:0] w3443;
	wire [0:0] w3444;
	wire [31:0] w3445;
	wire [0:0] w3447;
	wire [0:0] w3448;
	wire [31:0] w3449;
	wire [0:0] w3451;
	wire [0:0] w3452;
	wire [31:0] w3453;
	wire [0:0] w3455;
	wire [0:0] w3456;
	wire [31:0] w3457;
	wire [0:0] w3459;
	wire [31:0] w3460;
	wire [31:0] w3461;
	wire [0:0] w3462;
	wire [31:0] w3463;
	wire [31:0] w3464;
	wire [31:0] w3465;
	wire [31:0] w3466;
	wire [0:0] w3467;
	wire [31:0] w3468;
	wire [31:0] w3469;
	wire [31:0] w3470;
	wire [31:0] w3471;
	wire [31:0] w3472;
	wire [31:0] w3473;
	wire [31:0] w3474;
	wire [31:0] w3475;
	wire [0:0] w3476;
	wire [31:0] w3477;
	wire [31:0] w3478;
	wire [31:0] w3479;
	wire [31:0] w3480;
	wire [31:0] w3481;
	wire [31:0] w3482;
	wire [31:0] w3483;
	wire [31:0] w3484;
	wire [31:0] w3485;
	wire [31:0] w3486;
	wire [31:0] w3487;
	wire [31:0] w3488;
	wire [31:0] w3489;
	wire [31:0] w3490;
	wire [31:0] w3491;
	wire [31:0] w3492;
	wire [0:0] w3493;
	wire [31:0] w3494;
	wire [0:0] w3495;
	wire [31:0] w3496;
	wire [31:0] w3497;
	wire [31:0] w3499;
	wire [0:0] w3501;
	wire [0:0] w3502;
	wire [0:0] w3503;
	wire [0:0] w3504;
	wire [6:0] w3506;
	wire [6:0] w3507;
	wire [6:0] w3508;
	wire [6:0] w3510;
	wire [6:0] w3511;
	wire [6:0] w3512;
	wire [6:0] w3513;
	wire [6:0] w3514;
	wire [31:0] w3516;
	wire [31:0] w3517;
	wire [31:0] w3518;
	wire [31:0] w3520;
	wire [31:0] w3521;
	wire [0:0] w3523;
	wire [1:0] w3524;
	wire [1:0] w3525;
	wire [0:0] w3527;
	wire [0:0] w3528;
	wire [0:0] w3529;
	wire [0:0] w3531;
	wire [0:0] w3533;
	wire [0:0] w3534;
	wire [0:0] w3535;
	wire [0:0] w3536;
	wire [0:0] w3537;
	wire [0:0] w3538;
	wire [0:0] w3539;
	wire [0:0] w3540;
	wire [32:0] w3542;
	wire [32:0] w3543;
	wire [32:0] w3544;
	wire [32:0] w3545;
	wire [32:0] w3546;
	wire [31:0] w3548;
	wire [31:0] w3549;
	wire [31:0] w3550;
	wire [63:0] w3552;
	wire [63:0] w3553;
	wire [63:0] w3554;
	wire [63:0] w3556;
	wire [63:0] w3557;
	wire [63:0] w3558;
	wire [63:0] w3559;
	wire [63:0] w3561;
	wire [63:0] w3562;
	wire [6:0] w3563;
	wire [31:0] w3564;
	wire [0:0] w3565;
	wire [63:0] w3566;
	wire [63:0] w3567;
	wire [31:0] w3569;
	wire [31:0] w3570;
	wire [31:0] w3571;
	wire [31:0] w3572;
	wire [1:0] w3574;
	wire [4:0] w3576;
	wire [4:0] w3577;
	wire [4:0] w3578;
	wire [0:0] w3579;
	wire [0:0] w3580;
	wire [0:0] w3581;
	wire [4:0] w3582;
	wire [34:0] w3584;
	wire [33:0] w3586;
	wire [0:0] w3587;
	wire [34:0] w3588;
	wire [1:0] w3589;
	wire [0:0] w3590;
	wire [0:0] w3591;
	wire [0:0] w3592;
	wire [1:0] w3593;
	wire [0:0] w3594;
	wire [34:0] w3595;
	wire [16:0] w3596;
	wire [16:0] w3597;
	wire [16:0] w3598;
	wire [33:0] w3599;
	wire [0:0] w3600;
	wire [34:0] w3601;
	wire [0:0] w3602;
	wire [34:0] w3603;
	wire [16:0] w3604;
	wire [16:0] w3605;
	wire [33:0] w3606;
	wire [0:0] w3607;
	wire [34:0] w3608;
	wire [1:0] w3609;
	wire [0:0] w3610;
	wire [34:0] w3611;
	wire [34:0] w3612;
	wire [17:0] w3613;
	wire [15:0] w3614;
	wire [16:0] w3615;
	wire [34:0] w3616;
	wire [34:0] w3617;
	wire [34:0] w3618;
	wire [16:0] w3620;
	wire [16:0] w3621;
	wire [16:0] w3622;
	wire [1:0] w3624;
	wire [4:0] w3626;
	wire [4:0] w3627;
	wire [4:0] w3628;
	wire [0:0] w3629;
	wire [0:0] w3630;
	wire [4:0] w3631;
	wire [36:0] w3633;
	wire [35:0] w3635;
	wire [0:0] w3636;
	wire [36:0] w3637;
	wire [1:0] w3638;
	wire [0:0] w3639;
	wire [0:0] w3640;
	wire [0:0] w3641;
	wire [1:0] w3642;
	wire [0:0] w3643;
	wire [36:0] w3644;
	wire [17:0] w3645;
	wire [17:0] w3646;
	wire [17:0] w3647;
	wire [35:0] w3648;
	wire [0:0] w3649;
	wire [36:0] w3650;
	wire [0:0] w3651;
	wire [36:0] w3652;
	wire [17:0] w3653;
	wire [17:0] w3654;
	wire [35:0] w3655;
	wire [0:0] w3656;
	wire [36:0] w3657;
	wire [1:0] w3658;
	wire [0:0] w3659;
	wire [36:0] w3660;
	wire [36:0] w3661;
	wire [18:0] w3662;
	wire [17:0] w3663;
	wire [36:0] w3664;
	wire [36:0] w3665;
	wire [36:0] w3666;
	wire [17:0] w3668;
	wire [17:0] w3669;
	wire [1:0] w3671;
	wire [4:0] w3673;
	wire [4:0] w3674;
	wire [4:0] w3675;
	wire [0:0] w3676;
	wire [0:0] w3677;
	wire [4:0] w3678;
	wire [33:0] w3681;
	wire [0:0] w3682;
	wire [34:0] w3683;
	wire [1:0] w3684;
	wire [0:0] w3685;
	wire [0:0] w3686;
	wire [0:0] w3687;
	wire [1:0] w3688;
	wire [0:0] w3689;
	wire [34:0] w3690;
	wire [16:0] w3691;
	wire [16:0] w3692;
	wire [16:0] w3693;
	wire [33:0] w3694;
	wire [0:0] w3695;
	wire [34:0] w3696;
	wire [0:0] w3697;
	wire [34:0] w3698;
	wire [16:0] w3699;
	wire [16:0] w3700;
	wire [33:0] w3701;
	wire [0:0] w3702;
	wire [34:0] w3703;
	wire [1:0] w3704;
	wire [0:0] w3705;
	wire [34:0] w3706;
	wire [34:0] w3707;
	wire [15:0] w3708;
	wire [16:0] w3709;
	wire [34:0] w3710;
	wire [34:0] w3711;
	wire [34:0] w3712;
	wire [16:0] w3714;
	wire [16:0] w3715;
	wire [63:0] w3717;
	wire [63:0] w3718;
	wire [63:0] w3719;
	wire [63:0] w3720;
	wire [63:0] w3721;
	wire [31:0] w3724;
	wire [31:0] w3726;
	wire [7:0] w3728;
	wire [7:0] w3729;
	wire [7:0] w3731;
	wire [0:0] w3732;
	wire [0:0] w3733;
	wire [0:0] w3734;
	wire [0:0] w3735;
	wire [0:0] w3736;
	wire [0:0] w3737;
	wire [0:0] w3738;
	wire [0:0] w3739;
	wire [0:0] w3740;
	wire [0:0] w3741;
	wire [0:0] w3742;
	wire [0:0] w3743;
	wire [0:0] w3744;
	wire [0:0] w3745;
	wire [0:0] w3746;
	wire [0:0] w3747;
	wire [0:0] w3748;
	wire [0:0] w3749;
	wire [0:0] w3750;
	wire [0:0] w3751;
	wire [0:0] w3752;
	wire [0:0] w3753;
	wire [0:0] w3754;
	wire [0:0] w3755;
	wire [0:0] w3756;
	wire [0:0] w3757;
	wire [31:0] w3758;
	wire [0:0] w3760;
	wire [0:0] w3761;
	wire [0:0] w3762;
	wire [0:0] w3763;
	wire [0:0] w3764;
	wire [31:0] w3765;
	wire [0:0] w3768;
	wire [0:0] w3769;
	wire [0:0] w3770;
	wire [0:0] w3771;
	wire [0:0] w3772;
	wire [31:0] w3773;
	wire [0:0] w3775;
	wire [0:0] w3776;
	wire [0:0] w3777;
	wire [0:0] w3778;
	wire [31:0] w3779;
	wire [0:0] w3781;
	wire [0:0] w3782;
	wire [0:0] w3783;
	wire [0:0] w3784;
	wire [0:0] w3785;
	wire [31:0] w3786;
	wire [0:0] w3788;
	wire [0:0] w3789;
	wire [0:0] w3790;
	wire [31:0] w3791;
	wire [0:0] w3793;
	wire [0:0] w3794;
	wire [0:0] w3795;
	wire [31:0] w3796;
	wire [0:0] w3798;
	wire [0:0] w3799;
	wire [0:0] w3800;
	wire [31:0] w3801;
	wire [0:0] w3803;
	wire [0:0] w3804;
	wire [0:0] w3805;
	wire [0:0] w3806;
	wire [0:0] w3807;
	wire [31:0] w3808;
	wire [0:0] w3810;
	wire [0:0] w3811;
	wire [0:0] w3812;
	wire [31:0] w3813;
	wire [0:0] w3815;
	wire [0:0] w3816;
	wire [0:0] w3817;
	wire [31:0] w3818;
	wire [0:0] w3820;
	wire [0:0] w3821;
	wire [0:0] w3822;
	wire [31:0] w3823;
	wire [0:0] w3825;
	wire [0:0] w3826;
	wire [0:0] w3827;
	wire [0:0] w3828;
	wire [31:0] w3829;
	wire [0:0] w3831;
	wire [0:0] w3832;
	wire [0:0] w3833;
	wire [31:0] w3834;
	wire [0:0] w3836;
	wire [0:0] w3837;
	wire [0:0] w3838;
	wire [31:0] w3839;
	wire [0:0] w3841;
	wire [0:0] w3842;
	wire [0:0] w3843;
	wire [31:0] w3844;
	wire [0:0] w3846;
	wire [0:0] w3847;
	wire [0:0] w3848;
	wire [0:0] w3849;
	wire [0:0] w3850;
	wire [31:0] w3851;
	wire [0:0] w3853;
	wire [0:0] w3854;
	wire [31:0] w3855;
	wire [0:0] w3857;
	wire [0:0] w3858;
	wire [31:0] w3859;
	wire [0:0] w3861;
	wire [0:0] w3862;
	wire [31:0] w3863;
	wire [0:0] w3865;
	wire [0:0] w3866;
	wire [31:0] w3867;
	wire [0:0] w3869;
	wire [0:0] w3870;
	wire [31:0] w3871;
	wire [0:0] w3873;
	wire [0:0] w3874;
	wire [31:0] w3875;
	wire [0:0] w3877;
	wire [0:0] w3878;
	wire [31:0] w3879;
	wire [0:0] w3881;
	wire [0:0] w3882;
	wire [31:0] w3883;
	wire [0:0] w3885;
	wire [0:0] w3886;
	wire [31:0] w3887;
	wire [0:0] w3889;
	wire [0:0] w3890;
	wire [31:0] w3891;
	wire [0:0] w3893;
	wire [0:0] w3894;
	wire [31:0] w3895;
	wire [0:0] w3897;
	wire [0:0] w3898;
	wire [31:0] w3899;
	wire [0:0] w3901;
	wire [0:0] w3902;
	wire [31:0] w3903;
	wire [0:0] w3905;
	wire [0:0] w3906;
	wire [31:0] w3907;
	wire [0:0] w3909;
	wire [0:0] w3910;
	wire [31:0] w3911;
	wire [0:0] w3913;
	wire [0:0] w3914;
	wire [0:0] w3915;
	wire [0:0] w3916;
	wire [0:0] w3917;
	wire [31:0] w3918;
	wire [0:0] w3920;
	wire [0:0] w3921;
	wire [31:0] w3922;
	wire [0:0] w3924;
	wire [0:0] w3925;
	wire [31:0] w3926;
	wire [0:0] w3928;
	wire [0:0] w3929;
	wire [31:0] w3930;
	wire [0:0] w3932;
	wire [0:0] w3933;
	wire [31:0] w3934;
	wire [0:0] w3936;
	wire [0:0] w3937;
	wire [31:0] w3938;
	wire [0:0] w3940;
	wire [0:0] w3941;
	wire [31:0] w3942;
	wire [0:0] w3944;
	wire [0:0] w3945;
	wire [31:0] w3946;
	wire [0:0] w3948;
	wire [0:0] w3949;
	wire [31:0] w3950;
	wire [0:0] w3952;
	wire [0:0] w3953;
	wire [31:0] w3954;
	wire [0:0] w3956;
	wire [0:0] w3957;
	wire [31:0] w3958;
	wire [0:0] w3960;
	wire [0:0] w3961;
	wire [31:0] w3962;
	wire [0:0] w3964;
	wire [0:0] w3965;
	wire [31:0] w3966;
	wire [0:0] w3968;
	wire [0:0] w3969;
	wire [31:0] w3970;
	wire [0:0] w3972;
	wire [0:0] w3973;
	wire [31:0] w3974;
	wire [0:0] w3976;
	wire [0:0] w3977;
	wire [31:0] w3978;
	wire [0:0] w3980;
	wire [0:0] w3981;
	wire [0:0] w3982;
	wire [0:0] w3983;
	wire [31:0] w3984;
	wire [0:0] w3986;
	wire [0:0] w3987;
	wire [31:0] w3988;
	wire [0:0] w3990;
	wire [0:0] w3991;
	wire [31:0] w3992;
	wire [0:0] w3994;
	wire [0:0] w3995;
	wire [31:0] w3996;
	wire [0:0] w3998;
	wire [0:0] w3999;
	wire [31:0] w4000;
	wire [0:0] w4002;
	wire [0:0] w4003;
	wire [31:0] w4004;
	wire [0:0] w4006;
	wire [0:0] w4007;
	wire [31:0] w4008;
	wire [0:0] w4010;
	wire [0:0] w4011;
	wire [31:0] w4012;
	wire [0:0] w4014;
	wire [0:0] w4015;
	wire [31:0] w4016;
	wire [0:0] w4018;
	wire [0:0] w4019;
	wire [31:0] w4020;
	wire [0:0] w4022;
	wire [0:0] w4023;
	wire [31:0] w4024;
	wire [0:0] w4026;
	wire [0:0] w4027;
	wire [31:0] w4028;
	wire [0:0] w4030;
	wire [0:0] w4031;
	wire [31:0] w4032;
	wire [0:0] w4034;
	wire [0:0] w4035;
	wire [31:0] w4036;
	wire [0:0] w4038;
	wire [0:0] w4039;
	wire [31:0] w4040;
	wire [0:0] w4042;
	wire [0:0] w4043;
	wire [31:0] w4044;
	wire [0:0] w4046;
	wire [0:0] w4047;
	wire [0:0] w4048;
	wire [0:0] w4049;
	wire [0:0] w4050;
	wire [31:0] w4051;
	wire [0:0] w4053;
	wire [0:0] w4054;
	wire [31:0] w4055;
	wire [0:0] w4057;
	wire [0:0] w4058;
	wire [31:0] w4059;
	wire [0:0] w4061;
	wire [0:0] w4062;
	wire [31:0] w4063;
	wire [0:0] w4065;
	wire [0:0] w4066;
	wire [31:0] w4067;
	wire [0:0] w4069;
	wire [0:0] w4070;
	wire [31:0] w4071;
	wire [0:0] w4073;
	wire [0:0] w4074;
	wire [31:0] w4075;
	wire [0:0] w4077;
	wire [0:0] w4078;
	wire [31:0] w4079;
	wire [0:0] w4081;
	wire [0:0] w4082;
	wire [31:0] w4083;
	wire [0:0] w4085;
	wire [0:0] w4086;
	wire [31:0] w4087;
	wire [0:0] w4089;
	wire [0:0] w4090;
	wire [31:0] w4091;
	wire [0:0] w4093;
	wire [0:0] w4094;
	wire [31:0] w4095;
	wire [0:0] w4097;
	wire [0:0] w4098;
	wire [31:0] w4099;
	wire [0:0] w4101;
	wire [0:0] w4102;
	wire [31:0] w4103;
	wire [0:0] w4105;
	wire [0:0] w4106;
	wire [31:0] w4107;
	wire [0:0] w4109;
	wire [0:0] w4110;
	wire [31:0] w4111;
	wire [0:0] w4113;
	wire [0:0] w4114;
	wire [0:0] w4115;
	wire [31:0] w4116;
	wire [0:0] w4118;
	wire [0:0] w4119;
	wire [31:0] w4120;
	wire [0:0] w4122;
	wire [0:0] w4123;
	wire [31:0] w4124;
	wire [0:0] w4126;
	wire [0:0] w4127;
	wire [31:0] w4128;
	wire [0:0] w4130;
	wire [0:0] w4131;
	wire [31:0] w4132;
	wire [0:0] w4134;
	wire [0:0] w4135;
	wire [31:0] w4136;
	wire [0:0] w4138;
	wire [0:0] w4139;
	wire [31:0] w4140;
	wire [0:0] w4142;
	wire [0:0] w4143;
	wire [31:0] w4144;
	wire [0:0] w4146;
	wire [0:0] w4147;
	wire [31:0] w4148;
	wire [0:0] w4150;
	wire [0:0] w4151;
	wire [31:0] w4152;
	wire [0:0] w4154;
	wire [0:0] w4155;
	wire [31:0] w4156;
	wire [0:0] w4158;
	wire [0:0] w4159;
	wire [31:0] w4160;
	wire [0:0] w4162;
	wire [0:0] w4163;
	wire [31:0] w4164;
	wire [0:0] w4166;
	wire [0:0] w4167;
	wire [31:0] w4168;
	wire [0:0] w4170;
	wire [0:0] w4171;
	wire [31:0] w4172;
	wire [0:0] w4174;
	wire [0:0] w4175;
	wire [31:0] w4176;
	wire [0:0] w4178;
	wire [0:0] w4179;
	wire [0:0] w4180;
	wire [31:0] w4181;
	wire [0:0] w4183;
	wire [0:0] w4184;
	wire [31:0] w4185;
	wire [0:0] w4187;
	wire [0:0] w4188;
	wire [31:0] w4189;
	wire [0:0] w4191;
	wire [0:0] w4192;
	wire [31:0] w4193;
	wire [0:0] w4195;
	wire [0:0] w4196;
	wire [31:0] w4197;
	wire [0:0] w4199;
	wire [0:0] w4200;
	wire [31:0] w4201;
	wire [0:0] w4203;
	wire [0:0] w4204;
	wire [31:0] w4205;
	wire [0:0] w4207;
	wire [0:0] w4208;
	wire [31:0] w4209;
	wire [0:0] w4211;
	wire [0:0] w4212;
	wire [31:0] w4213;
	wire [0:0] w4215;
	wire [0:0] w4216;
	wire [31:0] w4217;
	wire [0:0] w4219;
	wire [0:0] w4220;
	wire [31:0] w4221;
	wire [0:0] w4223;
	wire [0:0] w4224;
	wire [31:0] w4225;
	wire [0:0] w4227;
	wire [0:0] w4228;
	wire [31:0] w4229;
	wire [0:0] w4231;
	wire [0:0] w4232;
	wire [31:0] w4233;
	wire [0:0] w4235;
	wire [0:0] w4236;
	wire [31:0] w4237;
	wire [0:0] w4239;
	wire [0:0] w4240;
	wire [31:0] w4241;
	wire [0:0] w4243;
	wire [0:0] w4244;
	wire [0:0] w4245;
	wire [31:0] w4246;
	wire [0:0] w4248;
	wire [0:0] w4249;
	wire [31:0] w4250;
	wire [0:0] w4252;
	wire [0:0] w4253;
	wire [31:0] w4254;
	wire [0:0] w4256;
	wire [0:0] w4257;
	wire [31:0] w4258;
	wire [0:0] w4260;
	wire [0:0] w4261;
	wire [31:0] w4262;
	wire [0:0] w4264;
	wire [0:0] w4265;
	wire [31:0] w4266;
	wire [0:0] w4268;
	wire [0:0] w4269;
	wire [31:0] w4270;
	wire [0:0] w4272;
	wire [0:0] w4273;
	wire [31:0] w4274;
	wire [0:0] w4276;
	wire [0:0] w4277;
	wire [31:0] w4278;
	wire [0:0] w4280;
	wire [0:0] w4281;
	wire [31:0] w4282;
	wire [0:0] w4284;
	wire [0:0] w4285;
	wire [31:0] w4286;
	wire [0:0] w4288;
	wire [0:0] w4289;
	wire [31:0] w4290;
	wire [0:0] w4292;
	wire [0:0] w4293;
	wire [31:0] w4294;
	wire [0:0] w4296;
	wire [0:0] w4297;
	wire [31:0] w4298;
	wire [0:0] w4300;
	wire [0:0] w4301;
	wire [31:0] w4302;
	wire [0:0] w4304;
	wire [0:0] w4305;
	wire [31:0] w4306;
	wire [0:0] w4308;
	wire [0:0] w4309;
	wire [0:0] w4310;
	wire [0:0] w4311;
	wire [0:0] w4312;
	wire [31:0] w4313;
	wire [0:0] w4315;
	wire [0:0] w4316;
	wire [31:0] w4317;
	wire [0:0] w4319;
	wire [0:0] w4320;
	wire [31:0] w4321;
	wire [0:0] w4323;
	wire [0:0] w4324;
	wire [31:0] w4325;
	wire [0:0] w4327;
	wire [0:0] w4328;
	wire [31:0] w4329;
	wire [0:0] w4331;
	wire [0:0] w4332;
	wire [31:0] w4333;
	wire [0:0] w4335;
	wire [0:0] w4336;
	wire [31:0] w4337;
	wire [0:0] w4339;
	wire [0:0] w4340;
	wire [31:0] w4341;
	wire [0:0] w4343;
	wire [0:0] w4344;
	wire [31:0] w4345;
	wire [0:0] w4347;
	wire [0:0] w4348;
	wire [31:0] w4349;
	wire [0:0] w4351;
	wire [0:0] w4352;
	wire [31:0] w4353;
	wire [0:0] w4355;
	wire [0:0] w4356;
	wire [31:0] w4357;
	wire [0:0] w4359;
	wire [0:0] w4360;
	wire [31:0] w4361;
	wire [0:0] w4363;
	wire [0:0] w4364;
	wire [31:0] w4365;
	wire [0:0] w4367;
	wire [0:0] w4368;
	wire [31:0] w4369;
	wire [0:0] w4371;
	wire [0:0] w4372;
	wire [31:0] w4373;
	wire [0:0] w4375;
	wire [0:0] w4376;
	wire [0:0] w4377;
	wire [31:0] w4378;
	wire [0:0] w4380;
	wire [0:0] w4381;
	wire [31:0] w4382;
	wire [0:0] w4384;
	wire [0:0] w4385;
	wire [31:0] w4386;
	wire [0:0] w4388;
	wire [0:0] w4389;
	wire [31:0] w4390;
	wire [0:0] w4392;
	wire [0:0] w4393;
	wire [31:0] w4394;
	wire [0:0] w4396;
	wire [0:0] w4397;
	wire [31:0] w4398;
	wire [0:0] w4400;
	wire [0:0] w4401;
	wire [31:0] w4402;
	wire [0:0] w4404;
	wire [0:0] w4405;
	wire [31:0] w4406;
	wire [0:0] w4408;
	wire [0:0] w4409;
	wire [31:0] w4410;
	wire [0:0] w4412;
	wire [0:0] w4413;
	wire [31:0] w4414;
	wire [0:0] w4416;
	wire [0:0] w4417;
	wire [31:0] w4418;
	wire [0:0] w4420;
	wire [0:0] w4421;
	wire [31:0] w4422;
	wire [0:0] w4424;
	wire [0:0] w4425;
	wire [31:0] w4426;
	wire [0:0] w4428;
	wire [0:0] w4429;
	wire [31:0] w4430;
	wire [0:0] w4432;
	wire [0:0] w4433;
	wire [31:0] w4434;
	wire [0:0] w4436;
	wire [0:0] w4437;
	wire [31:0] w4438;
	wire [0:0] w4440;
	wire [0:0] w4441;
	wire [0:0] w4442;
	wire [31:0] w4443;
	wire [0:0] w4445;
	wire [0:0] w4446;
	wire [31:0] w4447;
	wire [0:0] w4449;
	wire [0:0] w4450;
	wire [31:0] w4451;
	wire [0:0] w4453;
	wire [0:0] w4454;
	wire [31:0] w4455;
	wire [0:0] w4457;
	wire [0:0] w4458;
	wire [31:0] w4459;
	wire [0:0] w4461;
	wire [0:0] w4462;
	wire [31:0] w4463;
	wire [0:0] w4465;
	wire [0:0] w4466;
	wire [31:0] w4467;
	wire [0:0] w4469;
	wire [0:0] w4470;
	wire [31:0] w4471;
	wire [0:0] w4473;
	wire [0:0] w4474;
	wire [31:0] w4475;
	wire [0:0] w4477;
	wire [0:0] w4478;
	wire [31:0] w4479;
	wire [0:0] w4481;
	wire [0:0] w4482;
	wire [31:0] w4483;
	wire [0:0] w4485;
	wire [0:0] w4486;
	wire [31:0] w4487;
	wire [0:0] w4489;
	wire [0:0] w4490;
	wire [31:0] w4491;
	wire [0:0] w4493;
	wire [0:0] w4494;
	wire [31:0] w4495;
	wire [0:0] w4497;
	wire [0:0] w4498;
	wire [31:0] w4499;
	wire [0:0] w4501;
	wire [0:0] w4502;
	wire [31:0] w4503;
	wire [0:0] w4505;
	wire [0:0] w4506;
	wire [0:0] w4507;
	wire [31:0] w4508;
	wire [0:0] w4510;
	wire [0:0] w4511;
	wire [31:0] w4512;
	wire [0:0] w4514;
	wire [0:0] w4515;
	wire [31:0] w4516;
	wire [0:0] w4518;
	wire [0:0] w4519;
	wire [31:0] w4520;
	wire [0:0] w4522;
	wire [0:0] w4523;
	wire [31:0] w4524;
	wire [0:0] w4526;
	wire [0:0] w4527;
	wire [31:0] w4528;
	wire [0:0] w4530;
	wire [0:0] w4531;
	wire [31:0] w4532;
	wire [0:0] w4534;
	wire [0:0] w4535;
	wire [31:0] w4536;
	wire [0:0] w4538;
	wire [0:0] w4539;
	wire [31:0] w4540;
	wire [0:0] w4542;
	wire [0:0] w4543;
	wire [31:0] w4544;
	wire [0:0] w4546;
	wire [0:0] w4547;
	wire [31:0] w4548;
	wire [0:0] w4550;
	wire [0:0] w4551;
	wire [31:0] w4552;
	wire [0:0] w4554;
	wire [0:0] w4555;
	wire [31:0] w4556;
	wire [0:0] w4558;
	wire [0:0] w4559;
	wire [31:0] w4560;
	wire [0:0] w4562;
	wire [0:0] w4563;
	wire [31:0] w4564;
	wire [0:0] w4566;
	wire [0:0] w4567;
	wire [31:0] w4568;
	wire [0:0] w4570;
	wire [0:0] w4571;
	wire [0:0] w4572;
	wire [0:0] w4573;
	wire [31:0] w4574;
	wire [0:0] w4576;
	wire [0:0] w4577;
	wire [31:0] w4578;
	wire [0:0] w4580;
	wire [0:0] w4581;
	wire [31:0] w4582;
	wire [0:0] w4584;
	wire [0:0] w4585;
	wire [31:0] w4586;
	wire [0:0] w4588;
	wire [0:0] w4589;
	wire [31:0] w4590;
	wire [0:0] w4592;
	wire [0:0] w4593;
	wire [31:0] w4594;
	wire [0:0] w4596;
	wire [0:0] w4597;
	wire [31:0] w4598;
	wire [0:0] w4600;
	wire [0:0] w4601;
	wire [31:0] w4602;
	wire [0:0] w4604;
	wire [0:0] w4605;
	wire [31:0] w4606;
	wire [0:0] w4608;
	wire [0:0] w4609;
	wire [31:0] w4610;
	wire [0:0] w4612;
	wire [0:0] w4613;
	wire [31:0] w4614;
	wire [0:0] w4616;
	wire [0:0] w4617;
	wire [31:0] w4618;
	wire [0:0] w4620;
	wire [0:0] w4621;
	wire [31:0] w4622;
	wire [0:0] w4624;
	wire [0:0] w4625;
	wire [31:0] w4626;
	wire [0:0] w4628;
	wire [0:0] w4629;
	wire [31:0] w4630;
	wire [0:0] w4632;
	wire [0:0] w4633;
	wire [31:0] w4634;
	wire [0:0] w4636;
	wire [0:0] w4637;
	wire [0:0] w4638;
	wire [31:0] w4639;
	wire [0:0] w4641;
	wire [0:0] w4642;
	wire [31:0] w4643;
	wire [0:0] w4645;
	wire [0:0] w4646;
	wire [31:0] w4647;
	wire [0:0] w4649;
	wire [0:0] w4650;
	wire [31:0] w4651;
	wire [0:0] w4653;
	wire [0:0] w4654;
	wire [31:0] w4655;
	wire [0:0] w4657;
	wire [0:0] w4658;
	wire [31:0] w4659;
	wire [0:0] w4661;
	wire [0:0] w4662;
	wire [31:0] w4663;
	wire [0:0] w4665;
	wire [0:0] w4666;
	wire [31:0] w4667;
	wire [0:0] w4669;
	wire [0:0] w4670;
	wire [31:0] w4671;
	wire [0:0] w4673;
	wire [0:0] w4674;
	wire [31:0] w4675;
	wire [0:0] w4677;
	wire [0:0] w4678;
	wire [31:0] w4679;
	wire [0:0] w4681;
	wire [0:0] w4682;
	wire [31:0] w4683;
	wire [0:0] w4685;
	wire [0:0] w4686;
	wire [31:0] w4687;
	wire [0:0] w4689;
	wire [0:0] w4690;
	wire [31:0] w4691;
	wire [0:0] w4693;
	wire [0:0] w4694;
	wire [31:0] w4695;
	wire [0:0] w4697;
	wire [0:0] w4698;
	wire [31:0] w4699;
	wire [0:0] w4701;
	wire [0:0] w4702;
	wire [0:0] w4703;
	wire [31:0] w4704;
	wire [0:0] w4706;
	wire [0:0] w4707;
	wire [31:0] w4708;
	wire [0:0] w4710;
	wire [0:0] w4711;
	wire [31:0] w4712;
	wire [0:0] w4714;
	wire [0:0] w4715;
	wire [31:0] w4716;
	wire [0:0] w4718;
	wire [0:0] w4719;
	wire [31:0] w4720;
	wire [0:0] w4722;
	wire [0:0] w4723;
	wire [31:0] w4724;
	wire [0:0] w4726;
	wire [0:0] w4727;
	wire [31:0] w4728;
	wire [0:0] w4730;
	wire [0:0] w4731;
	wire [31:0] w4732;
	wire [0:0] w4734;
	wire [0:0] w4735;
	wire [31:0] w4736;
	wire [0:0] w4738;
	wire [0:0] w4739;
	wire [31:0] w4740;
	wire [0:0] w4742;
	wire [0:0] w4743;
	wire [31:0] w4744;
	wire [0:0] w4746;
	wire [0:0] w4747;
	wire [31:0] w4748;
	wire [0:0] w4750;
	wire [0:0] w4751;
	wire [31:0] w4752;
	wire [0:0] w4754;
	wire [0:0] w4755;
	wire [31:0] w4756;
	wire [0:0] w4758;
	wire [0:0] w4759;
	wire [31:0] w4760;
	wire [0:0] w4762;
	wire [0:0] w4763;
	wire [31:0] w4764;
	wire [0:0] w4766;
	wire [0:0] w4767;
	wire [0:0] w4768;
	wire [31:0] w4769;
	wire [0:0] w4771;
	wire [0:0] w4772;
	wire [31:0] w4773;
	wire [0:0] w4775;
	wire [0:0] w4776;
	wire [31:0] w4777;
	wire [0:0] w4779;
	wire [0:0] w4780;
	wire [31:0] w4781;
	wire [0:0] w4783;
	wire [0:0] w4784;
	wire [31:0] w4785;
	wire [0:0] w4787;
	wire [0:0] w4788;
	wire [31:0] w4789;
	wire [0:0] w4791;
	wire [0:0] w4792;
	wire [31:0] w4793;
	wire [0:0] w4795;
	wire [0:0] w4796;
	wire [31:0] w4797;
	wire [0:0] w4799;
	wire [0:0] w4800;
	wire [31:0] w4801;
	wire [0:0] w4803;
	wire [0:0] w4804;
	wire [31:0] w4805;
	wire [0:0] w4807;
	wire [0:0] w4808;
	wire [31:0] w4809;
	wire [0:0] w4811;
	wire [0:0] w4812;
	wire [31:0] w4813;
	wire [0:0] w4815;
	wire [0:0] w4816;
	wire [31:0] w4817;
	wire [0:0] w4819;
	wire [0:0] w4820;
	wire [31:0] w4821;
	wire [0:0] w4823;
	wire [0:0] w4824;
	wire [31:0] w4825;
	wire [0:0] w4827;
	wire [0:0] w4828;
	wire [31:0] w4829;
	wire [31:0] w4831;
	wire [31:0] w4832;
	wire [31:0] w4834;
	wire [31:0] w4835;
	wire [0:0] w4837;
	wire [0:0] w4838;
	wire [0:0] w4839;
	wire [0:0] w4841;
	wire [0:0] w4842;
	wire [31:0] w4844;
	wire [31:0] w4845;
	wire [0:0] w4846;
	wire [31:0] w4847;
	wire [0:0] w4848;
	wire [31:0] w4849;
	wire [31:0] w4850;
	wire [31:0] w4852;
	wire [31:0] w4853;
	wire [0:0] w4854;
	wire [0:0] w4855;
	wire [0:0] w4856;
	wire [0:0] w4857;
	wire [0:0] w4858;
	wire [0:0] w4859;
	wire [0:0] w4861;
	wire [0:0] w4862;
	wire [0:0] w4863;
	wire [0:0] w4865;
	wire [0:0] w4866;
	wire [0:0] w4867;
	wire [0:0] w4869;
	wire [0:0] w4870;
	wire [31:0] w4872;
	wire [31:0] w4873;
	wire [31:0] w4875;
	wire [31:0] w4876;
	wire [31:0] w4878;
	wire [31:0] w4879;
	wire [31:0] w4880;
	wire [31:0] w4881;
	wire [31:0] w4883;
	wire [31:0] w4884;
	wire [31:0] w4885;
	wire [0:0] w4887;
	wire [0:0] w4888;
	wire [0:0] w4890;
	wire [0:0] w4891;
	wire [31:0] w4893;
	wire [31:0] w4894;
	wire [1:0] w4896;
	wire [29:0] w4897;
	wire [31:0] w4898;
	wire [31:0] w4899;
	wire [3:0] w4901;
	wire [3:0] w4902;
	wire [2:0] w4903;
	wire [3:0] w4904;
	wire [3:0] w4905;
	wire [3:0] w4906;
	wire [3:0] w4907;
	wire [3:0] w4908;
	wire [3:0] w4909;
	wire [1:0] w4910;
	wire [1:0] w4911;
	wire [3:0] w4912;
	wire [3:0] w4913;
	wire [2:0] w4914;
	wire [2:0] w4915;
	wire [3:0] w4916;
	wire [3:0] w4917;
	wire [3:0] w4918;
	wire [3:0] w4919;
	wire [3:0] w4920;
	wire [3:0] w4921;
	wire [3:0] w4922;
	wire [3:0] w4923;
	wire [3:0] w4924;
	wire [3:0] w4925;
	wire [3:0] w4926;
	wire [3:0] w4927;
	wire [31:0] w4929;
	wire [31:0] w4930;
	wire [31:0] w4932;
	wire [31:0] w4933;
	wire [0:0] w4935;
	wire [4:0] w4937;
	wire [4:0] w4938;
	wire [4:0] w4939;
	wire [4:0] w4940;
	wire [4:0] w4941;
	wire [4:0] w4942;
	wire [4:0] w4943;
	wire [4:0] w4944;
	wire [4:0] w4945;
	wire [30:0] w4947;
	wire [31:0] w4948;
	wire [31:0] w4949;
	wire [27:0] w4950;
	wire [31:0] w4951;
	wire [31:0] w4952;
	wire [31:0] w4953;
	wire [31:0] w4954;
	wire [30:0] w4956;
	wire [30:0] w4957;
	wire [30:0] w4958;
	wire [27:0] w4959;
	wire [0:0] w4960;
	wire [28:0] w4961;
	wire [0:0] w4962;
	wire [29:0] w4963;
	wire [0:0] w4964;
	wire [30:0] w4965;
	wire [30:0] w4966;
	wire [0:0] w4967;
	wire [31:0] w4968;
	wire [31:0] w4969;
	wire [31:0] w4970;
	wire [30:0] w4972;
	wire [31:0] w4973;
	wire [31:0] w4974;
	wire [27:0] w4975;
	wire [31:0] w4976;
	wire [31:0] w4977;
	wire [31:0] w4978;
	wire [31:0] w4979;
	wire [31:0] w4981;
	wire [31:0] w4982;
	wire [31:0] w4984;
	wire [31:0] w4985;
	wire [0:0] w4987;
	wire [31:0] w4988;
	wire [0:0] w4990;
	wire [31:0] w4991;

	// array write assignment wires

	// assignments
	assign w4991 = {w2011, w4990};
	assign w4985 = i13 ? w4984 : w117;
	assign w4976 = {w4975, w696};
	assign w4975 = s3001[27:0];
	assign w4973 = {w4972, w47};
	assign w4968 = {w4967, w4966};
	assign w4967 = s3000[31:31];
	assign w4963 = {w4962, w4961};
	assign w4962 = s3000[31:31];
	assign w4961 = {w4960, w4959};
	assign w4956 = s3000[30:0];
	assign w4952 = w3243 ? w4951 : w4949;
	assign w4950 = s2999[31:4];
	assign w4949 = w3240 ? w4948 : s2999;
	assign w4942 = s2997 - w4941;
	assign w4941 = {2'b00, w44};
	assign w4939 = s2997 - w4938;
	assign w4938 = {4'b0000, w23};
	assign w4937 = w944[4:0];
	assign w4933 = i13 ? w4932 : w117;
	assign w4930 = i13 ? w4929 : w117;
	assign w4927 = i12 ? w4926 : s2760;
	assign w4926 = i13 ? w4925 : w696;
	assign w4923 = s55 ? w4922 : s2760;
	assign w4922 = w3187 ? w2577 : w4921;
	assign w4921 = w3184 ? w4918 : s2760;
	assign w4919 = w294 ? w4918 : s2760;
	assign w4917 = w3255 ? w4916 : w4913;
	assign w4916 = {w47, w4915};
	assign w4914 = 3'b010;
	assign w4912 = {w688, w4911};
	assign w4910 = w913 ? w688 : w32;
	assign w4909 = w3191 ? w4908 : w4905;
	assign w4908 = s55 ? w4907 : s2760;
	assign w4905 = w3177 ? w4904 : w4902;
	assign w4904 = {w47, w4903};
	assign w4902 = w3227 ? w4901 : s2760;
	assign w4899 = i13 ? w4898 : w117;
	assign w4898 = {w4897, w4896};
	assign w4896 = {s2702, s2700};
	assign w4890 = w2721 ? w47 : s2615;
	assign w4888 = i13 ? w4887 : w47;
	assign w4885 = i13 ? w4884 : w117;
	assign w4883 = s2729 | s2632;
	assign w4880 = w4854 ? w117 : w4879;
	assign w4876 = i13 ? w4875 : w117;
	assign w4873 = i13 ? w4872 : w117;
	assign w4870 = i13 ? w4869 : w47;
	assign w4867 = i13 ? w4866 : s2612;
	assign w4866 = s2601 ? w23 : w4865;
	assign w4862 = w4848 ? w4861 : s2611;
	assign w4856 = ~i13;
	assign w4853 = s2596 - w4852;
	assign w4852 = {31'b0000000000000000000000000000000, w23};
	assign w4850 = i13 ? w4849 : w117;
	assign w4846 = s2606 == s2617;
	assign w4842 = i13 ? w4841 : w47;
	assign w4841 = w2721 ? w23 : w47;
	assign w4925 = w982 ? w4924 : w4901;
	assign w4839 = i13 ? w4838 : w47;
	assign w4838 = s2601 ? w23 : w4837;
	assign w4837 = s2611 ? w47 : s2600;
	assign w4834 = w2721 ? s18 : w117;
	assign w4832 = i13 ? w4831 : w117;
	assign w4831 = s2600 ? s2597 : w117;
	assign w4829 = w4828 ? w3726 : s2001;
	assign w4827 = w3841 & w4766;
	assign w4821 = w4820 ? w3726 : s1998;
	assign w4812 = w4811 & w3756;
	assign w4809 = w4808 ? w3726 : s1993;
	assign w4807 = w3815 & w4766;
	assign w4805 = w4804 ? w3726 : s1991;
	assign w4804 = w4803 & w3756;
	assign w4799 = w3805 & w4766;
	assign w4792 = w4791 & w3756;
	assign w4789 = w4788 ? w3726 : s1983;
	assign w4788 = w4787 & w3756;
	assign w4787 = w3788 & w4766;
	assign w4785 = w4784 ? w3726 : s1982;
	assign w4784 = w4783 & w3756;
	assign w4776 = w4775 & w3756;
	assign w4775 = w3770 & w4766;
	assign w4769 = w4768 ? w3726 : s1975;
	assign w4767 = w3742 & w4766;
	assign w4766 = w3980 & w4570;
	assign w4763 = w4762 & w3756;
	assign w4760 = w4759 ? w3726 : s1969;
	assign w4754 = w3831 & w4701;
	assign w4752 = w4751 ? w3726 : s1966;
	assign w4751 = w4750 & w3756;
	assign w4748 = w4747 ? w3726 : s1963;
	assign w4747 = w4746 & w3756;
	assign w4780 = w4779 & w3756;
	assign w4742 = w3815 & w4701;
	assign w4740 = w4739 ? w3726 : s1960;
	assign w4739 = w4738 & w3756;
	assign w4736 = w4735 ? w3726 : s1959;
	assign w4735 = w4734 & w3756;
	assign w4734 = w3805 & w4701;
	assign w4732 = w4731 ? w3726 : s1955;
	assign w4731 = w4730 & w3756;
	assign w4728 = w4727 ? w3726 : s1954;
	assign w4726 = w3793 & w4701;
	assign w4724 = w4723 ? w3726 : s1952;
	assign w4723 = w4722 & w3756;
	assign w4722 = w3788 & w4701;
	assign w4718 = w3783 & w4701;
	assign w4712 = w4711 ? w3726 : s1947;
	assign w4707 = w4706 & w3756;
	assign w4701 = w3914 & w4570;
	assign w4698 = w4697 & w3756;
	assign w4695 = w4694 ? w3726 : s1937;
	assign w4693 = w3836 & w4636;
	assign w4690 = w4689 & w3756;
	assign w4689 = w3831 & w4636;
	assign w4686 = w4685 & w3756;
	assign w4683 = w4682 ? w3726 : s1931;
	assign w4681 = w3820 & w4636;
	assign w4679 = w4678 ? w3726 : s1930;
	assign w4678 = w4677 & w3756;
	assign w4674 = w4673 & w3756;
	assign w4673 = w3810 & w4636;
	assign w4671 = w4670 ? w3726 : s1927;
	assign w4667 = w4666 ? w3726 : s1923;
	assign w4666 = w4665 & w3756;
	assign w4663 = w4662 ? w3726 : s1922;
	assign w4661 = w3793 & w4636;
	assign w4659 = w4658 ? w3726 : s1920;
	assign w4658 = w4657 & w3756;
	assign w4655 = w4654 ? w3726 : s1919;
	assign w4819 = w3831 & w4766;
	assign w4649 = w3776 & w4636;
	assign w4647 = w4646 ? w3726 : s1915;
	assign w4801 = w4800 ? w3726 : s1990;
	assign w4645 = w3770 & w4636;
	assign w4643 = w4642 ? w3726 : s1913;
	assign w4641 = w3762 & w4636;
	assign w4638 = w4637 & w3756;
	assign w4633 = w4632 & w3756;
	assign w4632 = w3841 & w4571;
	assign w4630 = w4629 ? w3726 : s1906;
	assign w4628 = w3836 & w4571;
	assign w4626 = w4625 ? w3726 : s1904;
	assign w4625 = w4624 & w3756;
	assign w4622 = w4621 ? w3726 : s1903;
	assign w4621 = w4620 & w3756;
	assign w4620 = w3826 & w4571;
	assign w4618 = w4617 ? w3726 : s1900;
	assign w4617 = w4616 & w3756;
	assign w4911 = w2754 ? w34 : w4910;
	assign w4616 = w3820 & w4571;
	assign w4613 = w4612 & w3756;
	assign w4612 = w3815 & w4571;
	assign w4608 = w3810 & w4571;
	assign w4605 = w4604 & w3756;
	assign w4601 = w4600 & w3756;
	assign w4598 = w4597 ? w3726 : s1891;
	assign w4597 = w4596 & w3756;
	assign w4594 = w4593 ? w3726 : s1889;
	assign w4593 = w4592 & w3756;
	assign w4592 = w3788 & w4571;
	assign w4590 = w4589 ? w3726 : s1888;
	assign w4589 = w4588 & w3756;
	assign w4588 = w3783 & w4571;
	assign w4586 = w4585 ? w3726 : s1885;
	assign w4584 = w3776 & w4571;
	assign w4582 = w4581 ? w3726 : s1884;
	assign w4581 = w4580 & w3756;
	assign w4580 = w3770 & w4571;
	assign w4578 = w4577 ? w3726 : s1882;
	assign w4574 = w4573 ? w3726 : s1881;
	assign w4573 = w4572 & w3756;
	assign w4570 = w4046 & w4308;
	assign w4567 = w4566 & w3756;
	assign w4564 = w4563 ? w3726 : s1873;
	assign w4563 = w4562 & w3756;
	assign w4560 = w4559 ? w3726 : s1871;
	assign w4558 = w3831 & w4505;
	assign w4556 = w4555 ? w3726 : s1870;
	assign w4554 = w3826 & w4505;
	assign w4845 = s2606 + w4844;
	assign w4551 = w4550 & w3756;
	assign w4547 = w4546 & w3756;
	assign w4539 = w4538 & w3756;
	assign w4536 = w4535 ? w3726 : s1859;
	assign w4531 = w4530 & w3756;
	assign w4527 = w4526 & w3756;
	assign w4524 = w4523 ? w3726 : s1855;
	assign w4522 = w3783 & w4505;
	assign w4520 = w4519 ? w3726 : s1852;
	assign w4516 = w4515 ? w3726 : s1851;
	assign w4514 = w3770 & w4505;
	assign w4506 = w3742 & w4505;
	assign w4505 = w3980 & w4309;
	assign w4501 = w3841 & w4440;
	assign w4499 = w4498 ? w3726 : s1842;
	assign w4495 = w4494 ? w3726 : s1840;
	assign w4530 = w3793 & w4505;
	assign w4486 = w4485 & w3756;
	assign w4483 = w4482 ? w3726 : s1835;
	assign w4482 = w4481 & w3756;
	assign w4479 = w4478 ? w3726 : s1833;
	assign w4478 = w4477 & w3756;
	assign w4477 = w3810 & w4440;
	assign w4783 = w3783 & w4766;
	assign w4475 = w4474 ? w3726 : s1832;
	assign w4474 = w4473 & w3756;
	assign w4465 = w3793 & w4440;
	assign w4463 = w4462 ? w3726 : s1825;
	assign w4462 = w4461 & w3756;
	assign w4461 = w3788 & w4440;
	assign w4459 = w4458 ? w3726 : s1824;
	assign w4458 = w4457 & w3756;
	assign w4457 = w3783 & w4440;
	assign w4510 = w3762 & w4505;
	assign w4455 = w4454 ? w3726 : s1821;
	assign w4614 = w4613 ? w3726 : s1899;
	assign w4451 = w4450 ? w3726 : s1820;
	assign w4447 = w4446 ? w3726 : s1818;
	assign w4446 = w4445 & w3756;
	assign w4443 = w4442 ? w3726 : s1817;
	assign w4442 = w4441 & w3756;
	assign w4438 = w4437 ? w3726 : s1811;
	assign w4437 = w4436 & w3756;
	assign w4436 = w3841 & w4375;
	assign w4434 = w4433 ? w3726 : s1810;
	assign w4432 = w3836 & w4375;
	assign w4429 = w4428 & w3756;
	assign w4424 = w3826 & w4375;
	assign w4422 = w4421 ? w3726 : s1804;
	assign w4414 = w4413 ? w3726 : s1801;
	assign w4412 = w3810 & w4375;
	assign w4409 = w4408 & w3756;
	assign w4406 = w4405 ? w3726 : s1796;
	assign w4858 = w4856 | w4857;
	assign w4405 = w4404 & w3756;
	assign w4401 = w4400 & w3756;
	assign w4400 = w3793 & w4375;
	assign w4398 = w4397 ? w3726 : s1793;
	assign w4396 = w3788 & w4375;
	assign w4394 = w4393 ? w3726 : s1792;
	assign w4388 = w3776 & w4375;
	assign w4385 = w4384 & w3756;
	assign w4559 = w4558 & w3756;
	assign w4382 = w4381 ? w3726 : s1786;
	assign w4381 = w4380 & w3756;
	assign w4378 = w4377 ? w3726 : s1785;
	assign w4377 = w4376 & w3756;
	assign w4369 = w4368 ? w3726 : s1779;
	assign w4368 = w4367 & w3756;
	assign w4365 = w4364 ? w3726 : s1777;
	assign w4360 = w4359 & w3756;
	assign w4356 = w4355 & w3756;
	assign w4353 = w4352 ? w3726 : s1772;
	assign w4352 = w4351 & w3756;
	assign w4347 = w3810 & w4310;
	assign w4384 = w3770 & w4375;
	assign w4337 = w4336 ? w3726 : s1764;
	assign w4336 = w4335 & w3756;
	assign w4335 = w3793 & w4310;
	assign w4333 = w4332 ? w3726 : s1762;
	assign w4332 = w4331 & w3756;
	assign w4331 = w3788 & w4310;
	assign w4328 = w4327 & w3756;
	assign w4325 = w4324 ? w3726 : s1758;
	assign w4321 = w4320 ? w3726 : s1757;
	assign w4320 = w4319 & w3756;
	assign w4317 = w4316 ? w3726 : s1755;
	assign w4316 = w4315 & w3756;
	assign w4312 = w4311 & w3756;
	assign w4308 = w3750 == w23;
	assign w4306 = w4305 ? w3726 : s1745;
	assign w4300 = w3836 & w4243;
	assign w4297 = w4296 & w3756;
	assign w4296 = w3831 & w4243;
	assign w4293 = w4292 & w3756;
	assign w4292 = w3826 & w4243;
	assign w4756 = w4755 ? w3726 : s1967;
	assign w4290 = w4289 ? w3726 : s1738;
	assign w4289 = w4288 & w3756;
	assign w4286 = w4285 ? w3726 : s1737;
	assign w4284 = w3815 & w4243;
	assign w4697 = w3841 & w4636;
	assign w4282 = w4281 ? w3726 : s1735;
	assign w4280 = w3810 & w4243;
	assign w4278 = w4277 ? w3726 : s1734;
	assign w4699 = w4698 ? w3726 : s1938;
	assign w4453 = w3776 & w4440;
	assign w4276 = w3805 & w4243;
	assign w4273 = w4272 & w3756;
	assign w4270 = w4269 ? w3726 : s1729;
	assign w4268 = w3793 & w4243;
	assign w4265 = w4264 & w3756;
	assign w4262 = w4261 ? w3726 : s1726;
	assign w4261 = w4260 & w3756;
	assign w4857 = ~s2600;
	assign w4260 = w3783 & w4243;
	assign w4258 = w4257 ? w3726 : s1723;
	assign w4254 = w4253 ? w3726 : s1722;
	assign w4249 = w4248 & w3756;
	assign w4241 = w4240 ? w3726 : s1714;
	assign w4240 = w4239 & w3756;
	assign w4239 = w3841 & w4178;
	assign w4236 = w4235 & w3756;
	assign w4232 = w4231 & w3756;
	assign w4231 = w3831 & w4178;
	assign w4229 = w4228 ? w3726 : s1710;
	assign w4228 = w4227 & w3756;
	assign w4224 = w4223 & w3756;
	assign w4223 = w3820 & w4178;
	assign w4221 = w4220 ? w3726 : s1706;
	assign w4220 = w4219 & w3756;
	assign w4217 = w4216 ? w3726 : s1704;
	assign w4243 = w3980 & w4047;
	assign w4213 = w4212 ? w3726 : s1703;
	assign w4367 = w3836 & w4310;
	assign w4211 = w3805 & w4178;
	assign w4209 = w4208 ? w3726 : s1699;
	assign w4523 = w4522 & w3756;
	assign w4208 = w4207 & w3756;
	assign w4207 = w3798 & w4178;
	assign w4204 = w4203 & w3756;
	assign w4201 = w4200 ? w3726 : s1696;
	assign w4526 = w3788 & w4505;
	assign w4199 = w3788 & w4178;
	assign w4197 = w4196 ? w3726 : s1695;
	assign w4195 = w3783 & w4178;
	assign w4824 = w4823 & w3756;
	assign w4188 = w4187 & w3756;
	assign w4988 = {w2011, w4987};
	assign w4185 = w4184 ? w3726 : s1689;
	assign w4184 = w4183 & w3756;
	assign w4183 = w3762 & w4178;
	assign w4585 = w4584 & w3756;
	assign w4181 = w4180 ? w3726 : s1688;
	assign w4179 = w3742 & w4178;
	assign w4175 = w4174 & w3756;
	assign w4174 = w3841 & w4113;
	assign w4795 = w3798 & w4766;
	assign w4172 = w4171 ? w3726 : s1681;
	assign w4171 = w4170 & w3756;
	assign w4170 = w3836 & w4113;
	assign w4168 = w4167 ? w3726 : s1679;
	assign w4167 = w4166 & w3756;
	assign w4163 = w4162 & w3756;
	assign w4160 = w4159 ? w3726 : s1675;
	assign w4159 = w4158 & w3756;
	assign w4158 = w3820 & w4113;
	assign w4155 = w4154 & w3756;
	assign w4154 = w3815 & w4113;
	assign w4152 = w4151 ? w3726 : s1672;
	assign w4854 = s2626 == w4853;
	assign w4151 = w4150 & w3756;
	assign w4150 = w3810 & w4113;
	assign w4148 = w4147 ? w3726 : s1671;
	assign w4515 = w4514 & w3756;
	assign w4147 = w4146 & w3756;
	assign w4146 = w3805 & w4113;
	assign w4144 = w4143 ? w3726 : s1667;
	assign w4143 = w4142 & w3756;
	assign w4140 = w4139 ? w3726 : s1666;
	assign w4139 = w4138 & w3756;
	assign w4135 = w4134 & w3756;
	assign w4130 = w3783 & w4113;
	assign w4128 = w4127 ? w3726 : s1660;
	assign w4123 = w4122 & w3756;
	assign w4116 = w4115 ? w3726 : s1656;
	assign w4714 = w3776 & w4701;
	assign w4115 = w4114 & w3756;
	assign w4113 = w3847 & w4047;
	assign w4110 = w4109 & w3756;
	assign w4650 = w4649 & w3756;
	assign w4107 = w4106 ? w3726 : s1650;
	assign w4106 = w4105 & w3756;
	assign w4105 = w3836 & w4048;
	assign w4408 = w3805 & w4375;
	assign w4101 = w3831 & w4048;
	assign w4091 = w4090 ? w3726 : s1643;
	assign w4089 = w3815 & w4048;
	assign w4087 = w4086 ? w3726 : s1641;
	assign w4083 = w4082 ? w3726 : s1640;
	assign w4082 = w4081 & w3756;
	assign w4081 = w3805 & w4048;
	assign w4421 = w4420 & w3756;
	assign w4078 = w4077 & w3756;
	assign w4077 = w3798 & w4048;
	assign w4073 = w3793 & w4048;
	assign w4071 = w4070 ? w3726 : s1633;
	assign w4069 = w3788 & w4048;
	assign w4067 = w4066 ? w3726 : s1632;
	assign w4066 = w4065 & w3756;
	assign w4187 = w3770 & w4178;
	assign w4065 = w3783 & w4048;
	assign w4063 = w4062 ? w3726 : s1629;
	assign w4062 = w4061 & w3756;
	assign w4059 = w4058 ? w3726 : s1628;
	assign w4058 = w4057 & w3756;
	assign w4355 = w3820 & w4310;
	assign w4055 = w4054 ? w3726 : s1626;
	assign w4054 = w4053 & w3756;
	assign w4051 = w4050 ? w3726 : s1625;
	assign w4049 = w3742 & w4048;
	assign w4269 = w4268 & w3756;
	assign w4048 = w3747 & w4047;
	assign w4047 = w4046 & w3751;
	assign w4044 = w4043 ? w3726 : s1617;
	assign w4043 = w4042 & w3756;
	assign w4111 = w4110 ? w3726 : s1651;
	assign w4040 = w4039 ? w3726 : s1616;
	assign w4036 = w4035 ? w3726 : s1614;
	assign w4032 = w4031 ? w3726 : s1613;
	assign w4687 = w4686 ? w3726 : s1934;
	assign w4026 = w3820 & w3981;
	assign w4022 = w3815 & w3981;
	assign w4020 = w4019 ? w3726 : s1607;
	assign w4018 = w3810 & w3981;
	assign w4016 = w4015 ? w3726 : s1606;
	assign w4012 = w4011 ? w3726 : s1602;
	assign w4006 = w3793 & w3981;
	assign w4467 = w4466 ? w3726 : s1827;
	assign w4004 = w4003 ? w3726 : s1599;
	assign w4003 = w4002 & w3756;
	assign w4000 = w3999 ? w3726 : s1598;
	assign w3998 = w3783 & w3981;
	assign w3992 = w3991 ? w3726 : s1594;
	assign w4413 = w4412 & w3756;
	assign w3990 = w3770 & w3981;
	assign w3988 = w3987 ? w3726 : s1592;
	assign w4235 = w3836 & w4178;
	assign w3987 = w3986 & w3756;
	assign w4319 = w3770 & w4310;
	assign w4118 = w3762 & w4113;
	assign w3986 = w3762 & w3981;
	assign w3983 = w3982 & w3756;
	assign w3980 = w3846 & w3913;
	assign w3978 = w3977 ? w3726 : s1586;
	assign w3977 = w3976 & w3756;
	assign w3972 = w3836 & w3915;
	assign w3970 = w3969 ? w3726 : s1583;
	assign w4768 = w4767 & w3756;
	assign w3969 = w3968 & w3756;
	assign w3968 = w3831 & w3915;
	assign w4817 = w4816 ? w3726 : s1997;
	assign w3964 = w3826 & w3915;
	assign w4669 = w3805 & w4636;
	assign w3962 = w3961 ? w3726 : s1579;
	assign w3961 = w3960 & w3756;
	assign w3960 = w3820 & w3915;
	assign w3958 = w3957 ? w3726 : s1578;
	assign w3957 = w3956 & w3756;
	assign w3956 = w3815 & w3915;
	assign w3954 = w3953 ? w3726 : s1576;
	assign w4746 = w3820 & w4701;
	assign w3952 = w3810 & w3915;
	assign w3950 = w3949 ? w3726 : s1575;
	assign w4893 = w2718 ? s2632 : s2705;
	assign w4191 = w3776 & w4178;
	assign w3948 = w3805 & w3915;
	assign w3944 = w3798 & w3915;
	assign w4657 = w3788 & w4636;
	assign w3942 = w3941 ? w3726 : s1570;
	assign w3938 = w3937 ? w3726 : s1568;
	assign w3937 = w3936 & w3756;
	assign w4445 = w3762 & w4440;
	assign w3930 = w3929 ? w3726 : s1564;
	assign w3929 = w3928 & w3756;
	assign w4875 = w2721 ? s762 : w117;
	assign w4600 = w3798 & w4571;
	assign w3928 = w3776 & w3915;
	assign w3926 = w3925 ? w3726 : s1563;
	assign w3925 = w3924 & w3756;
	assign w3924 = w3770 & w3915;
	assign w3922 = w3921 ? w3726 : s1561;
	assign w3921 = w3920 & w3756;
	assign w3917 = w3916 & w3756;
	assign w3916 = w3742 & w3915;
	assign w3915 = w3914 & w3752;
	assign w3911 = w3910 ? w3726 : s1553;
	assign w3910 = w3909 & w3756;
	assign w3909 = w3841 & w3848;
	assign w3901 = w3831 & w3848;
	assign w3899 = w3898 ? w3726 : s1549;
	assign w3898 = w3897 & w3756;
	assign w3897 = w3826 & w3848;
	assign w3895 = w3894 ? w3726 : s1546;
	assign w3894 = w3893 & w3756;
	assign w3891 = w3890 ? w3726 : s1545;
	assign w3966 = w3965 ? w3726 : s1582;
	assign w3887 = w3886 ? w3726 : s1543;
	assign w3883 = w3882 ? w3726 : s1542;
	assign w3882 = w3881 & w3756;
	assign w3881 = w3805 & w3848;
	assign w3879 = w3878 ? w3726 : s1538;
	assign w3877 = w3798 & w3848;
	assign w3874 = w3873 & w3756;
	assign w3865 = w3783 & w3848;
	assign w3861 = w3776 & w3848;
	assign w3859 = w3858 ? w3726 : s1530;
	assign w3858 = w3857 & w3756;
	assign w3857 = w3770 & w3848;
	assign w3854 = w3853 & w3756;
	assign w3851 = w3850 ? w3726 : s1527;
	assign w3850 = w3849 & w3756;
	assign w3849 = w3742 & w3848;
	assign w3847 = w3846 & w3746;
	assign w3846 = w3743 == w23;
	assign w3844 = w3843 ? w3726 : s1521;
	assign w3843 = w3842 & w3756;
	assign w4502 = w4501 & w3756;
	assign w3842 = w3841 & w3753;
	assign w3841 = w3775 & w3825;
	assign w3837 = w3836 & w3753;
	assign w3834 = w3833 ? w3726 : s1518;
	assign w3833 = w3832 & w3756;
	assign w3831 = w3761 & w3825;
	assign w3829 = w3828 ? w3726 : s1517;
	assign w3828 = w3827 & w3756;
	assign w3827 = w3826 & w3753;
	assign w3826 = w3736 & w3825;
	assign w3825 = w3781 & w3803;
	assign w3821 = w3820 & w3753;
	assign w3914 = w3744 & w3913;
	assign w3820 = w3775 & w3804;
	assign w3818 = w3817 ? w3726 : s1513;
	assign w3817 = w3816 & w3756;
	assign w3813 = w3812 ? w3726 : s1511;
	assign w3812 = w3811 & w3756;
	assign w3811 = w3810 & w3753;
	assign w3804 = w3738 & w3803;
	assign w3801 = w3800 ? w3726 : s1505;
	assign w4309 = w3749 & w4308;
	assign w3799 = w3798 & w3753;
	assign w3798 = w3775 & w3782;
	assign w3793 = w3769 & w3782;
	assign w3790 = w3789 & w3756;
	assign w3789 = w3788 & w3753;
	assign w3788 = w3761 & w3782;
	assign w3786 = w3785 ? w3726 : s1501;
	assign w3782 = w3781 & w3740;
	assign w3777 = w3776 & w3753;
	assign w3775 = w3760 & w3768;
	assign w3771 = w3770 & w3753;
	assign w4127 = w4126 & w3756;
	assign w3770 = w3769 & w3741;
	assign w3764 = w3763 & w3756;
	assign w4136 = w4135 ? w3726 : s1664;
	assign w3762 = w3761 & w3741;
	assign w3761 = w3760 & w3735;
	assign w3760 = w3732 == w23;
	assign w3757 = w3754 & w3756;
	assign w3751 = w3750 == w47;
	assign w3747 = w3744 & w3746;
	assign w4606 = w4605 ? w3726 : s1896;
	assign w3746 = w3745 == w47;
	assign w4759 = w4758 & w3756;
	assign w3745 = w3731[5:5];
	assign w3742 = w3736 & w3741;
	assign w3741 = w3738 & w3740;
	assign w3740 = w3739 == w47;
	assign w3739 = w3731[3:3];
	assign w4311 = w3742 & w4310;
	assign w3738 = w3737 == w47;
	assign w3736 = w3733 & w3735;
	assign w3734 = w3731[1:1];
	assign w3733 = w3732 == w47;
	assign w3731 = w775 ? i48 : w3729;
	assign w3726 = w775 ? i46 : w3724;
	assign w3718 = {63'b000000000000000000000000000000000000000000000000000000000000000, w23};
	assign w3714 = w1310 ? w1303 : s1305;
	assign w3712 = i13 ? w3711 : w3584;
	assign w3704 = {1'b0, w23};
	assign w3946 = w3945 ? w3726 : s1571;
	assign w3701 = {w3699, w3700};
	assign w3699 = w3691 + s1305;
	assign w3698 = w3697 ? w3696 : w3690;
	assign w3697 = w3684 == w32;
	assign w3696 = {w3695, w3694};
	assign w4178 = w3914 & w4047;
	assign w3695 = w3692[16:16];
	assign w3693 = s1294[17:1];
	assign w3689 = |w3688;
	assign w3686 = |w3684;
	assign w3685 = w3684 == w34;
	assign w3683 = {w3682, w3681};
	assign w3675 = w1312 ? w3674 : s1270;
	assign w3673 = {4'b0000, w23};
	assign w4848 = s2609 & s2600;
	assign w3671 = i13 ? w1283 : w688;
	assign w3668 = w1259 ? w1252 : s1254;
	assign w3664 = {w3662, w3663};
	assign w3661 = w1261 ? w3660 : s1234;
	assign w3659 = w3638 == w3658;
	assign w3658 = {1'b0, w23};
	assign w4637 = w3742 & w4636;
	assign w3657 = {w3656, w3655};
	assign w3655 = {w3653, w3654};
	assign w3653 = w3645 + s1254;
	assign w3652 = w3651 ? w3650 : w3644;
	assign w3651 = w3638 == w32;
	assign w3677 = w3579 | w3676;
	assign w3650 = {w3649, w3648};
	assign w4665 = w3798 & w4636;
	assign w3649 = w3646[17:17];
	assign w3646 = w3645 + w1257;
	assign w3769 = w3733 & w3768;
	assign w3645 = s1234[36:19];
	assign w3644 = w3643 ? w3637 : i43;
	assign w3643 = |w3642;
	assign w3642 = {w3641, w3639};
	assign w4203 = w3793 & w4178;
	assign w3640 = |w3638;
	assign w3638 = s1234[1:0];
	assign w3635 = s1234[36:1];
	assign w3633 = 37'b0000000000000000000000000000000000000;
	assign w3627 = s1207 + w3626;
	assign w3626 = {4'b0000, w23};
	assign w4392 = w3783 & w4375;
	assign w3617 = w1196 ? w3616 : w3612;
	assign w4552 = w4551 ? w3726 : s1867;
	assign w3616 = {w3613, w3615};
	assign w3615 = {w3614, w47};
	assign w3613 = 18'b000000000000000000;
	assign w3886 = w3885 & w3756;
	assign w3611 = w3610 ? w3608 : w3603;
	assign w3609 = {1'b0, w23};
	assign w3606 = {w3604, w3605};
	assign w3605 = s1160[17:1];
	assign w3604 = w3596 + s1191;
	assign w3603 = w3602 ? w3601 : w3595;
	assign w3601 = {w3600, w3599};
	assign w3597 = w3596 + w1194;
	assign w3596 = s1160[34:18];
	assign w3593 = {w3592, w3590};
	assign w3592 = ~w3591;
	assign w3588 = {w3587, w3586};
	assign w3587 = s1160[34:34];
	assign w3584 = 35'b00000000000000000000000000000000000;
	assign w4543 = w4542 & w3756;
	assign w3581 = w3579 | w3580;
	assign w3578 = w1198 ? w3577 : s1134;
	assign w3577 = s1134 + w3576;
	assign w3595 = w3594 ? w3588 : i42;
	assign w3574 = i13 ? w1147 : w688;
	assign w3572 = i13 ? w3571 : w117;
	assign w3571 = w3565 ? w117 : w3570;
	assign w3570 = s1069 + w3569;
	assign w3567 = i13 ? w3566 : w1042;
	assign w3565 = s1069 == w3564;
	assign w4629 = w4628 & w3756;
	assign w3564 = {25'b0000000000000000000000000, w3563};
	assign w3563 = 7'b1100100;
	assign w3562 = s1043 + w3561;
	assign w4327 = w3783 & w4310;
	assign w3557 = s1011 + w3556;
	assign w3556 = {63'b000000000000000000000000000000000000000000000000000000000000000, w23};
	assign w3554 = i13 ? w3553 : w1042;
	assign w3550 = i13 ? w3549 : w117;
	assign w3784 = w3783 & w3753;
	assign w3545 = w3543 + w3544;
	assign w3544 = {1'b0, w944};
	assign w3542 = 33'b000000000000000000000000000000000;
	assign w3536 = w2746 ? s900 : w23;
	assign w3534 = w2754 ? w47 : w3533;
	assign w3533 = w913 ? w47 : s900;
	assign w3531 = i13 ? s900 : w47;
	assign w3779 = w3778 ? w3726 : s1497;
	assign w3529 = i13 ? w3528 : w47;
	assign w4471 = w4470 ? w3726 : s1828;
	assign w3524 = {w3523, w884};
	assign w3523 = s885[0:0];
	assign w3521 = i13 ? w3520 : w117;
	assign w3768 = w3734 == w23;
	assign w3518 = i13 ? w3517 : w117;
	assign w3514 = w775 ? w791 : w3513;
	assign w3513 = w802 ? s797 : w3512;
	assign w3512 = w808 ? w3511 : s797;
	assign w4466 = w4465 & w3756;
	assign w3511 = s797 + w3510;
	assign w3510 = {6'b000000, w23};
	assign w3641 = ~w3640;
	assign w3507 = w802 ? w3506 : s792;
	assign w3589 = s1160[1:0];
	assign w3506 = w796[6:0];
	assign w4277 = w4276 & w3756;
	assign w3504 = i12 ? w3503 : w47;
	assign w3503 = i13 ? w3502 : s772;
	assign w3501 = w3195 ? w811 : s772;
	assign w3495 = |w760;
	assign w3853 = w3762 & w3848;
	assign w3494 = w3493 ? w3492 : w3477;
	assign w3487 = w3462 ? w3486 : w3485;
	assign w3483 = w3462 ? w3482 : w3481;
	assign w3481 = w3459 ? s458 : s457;
	assign w3480 = w3462 ? w3479 : w3478;
	assign w4402 = w4401 ? w3726 : s1795;
	assign w3479 = w3459 ? s456 : s455;
	assign w4176 = w4175 ? w3726 : s1682;
	assign w3477 = w3476 ? w3475 : w3468;
	assign w3476 = w760[3:3];
	assign w3475 = w3467 ? w3474 : w3471;
	assign w3472 = w3459 ? s442 : s441;
	assign w3470 = w3459 ? s440 : s439;
	assign w3469 = w3459 ? s438 : s437;
	assign w3466 = w3462 ? w3465 : w3464;
	assign w3464 = w3459 ? s420 : s419;
	assign w3463 = w3462 ? w3461 : w3460;
	assign w3462 = w760[1:1];
	assign w3460 = w3459 ? s416 : s415;
	assign w3459 = w760[0:0];
	assign w3457 = w3456 ? w3293 : s475;
	assign w3455 = w3329 & w3442;
	assign w4793 = w4792 ? w3726 : s1985;
	assign w3452 = w3451 & w3313;
	assign w3449 = w3448 ? w3293 : s473;
	assign w3448 = w3447 & w3313;
	assign w3439 = w3438 & w3313;
	assign w3436 = w3435 ? w3293 : s470;
	assign w3435 = w3434 & w3313;
	assign w3434 = w3324 & w3425;
	assign w3965 = w3964 & w3756;
	assign w3432 = w3431 ? w3293 : s469;
	assign w3430 = w3318 & w3425;
	assign w3428 = w3427 ? w3293 : s468;
	assign w4924 = w3195 ? w4923 : w4920;
	assign w4248 = w3762 & w4243;
	assign w3427 = w3426 & w3313;
	assign w3422 = w3421 ? w3293 : s460;
	assign w3421 = w3420 & w3313;
	assign w4237 = w4236 ? w3726 : s1713;
	assign w3418 = w3417 ? w3293 : s459;
	assign w3416 = w3324 & w3407;
	assign w3413 = w3412 & w3313;
	assign w3407 = w3334 & w3389;
	assign w3405 = w3404 ? w3293 : s456;
	assign w3404 = w3403 & w3313;
	assign w3403 = w3329 & w3390;
	assign w3400 = w3399 & w3313;
	assign w3397 = w3396 ? w3293 : s454;
	assign w3390 = w3304 & w3389;
	assign w3389 = w3306 & w3388;
	assign w3388 = w3307 == w23;
	assign w3386 = w3385 ? w3293 : s444;
	assign w3385 = w3384 & w3313;
	assign w3489 = w3459 ? s475 : s474;
	assign w3382 = w3381 ? w3293 : s443;
	assign w3913 = w3745 == w23;
	assign w3381 = w3380 & w3313;
	assign w3380 = w3324 & w3371;
	assign w3376 = w3318 & w3371;
	assign w3373 = w3372 & w3313;
	assign w3369 = w3368 ? w3293 : s440;
	assign w3368 = w3367 & w3313;
	assign w3365 = w3364 ? w3293 : s439;
	assign w3363 = w3324 & w3354;
	assign w3357 = w3356 ? w3293 : s437;
	assign w3355 = w3302 & w3354;
	assign w3354 = w3304 & w3353;
	assign w4716 = w4715 ? w3726 : s1948;
	assign w3543 = {1'b0, s18};
	assign w3353 = w3352 & w3308;
	assign w3352 = w3305 == w23;
	assign w3350 = w3349 ? w3293 : s422;
	assign w3348 = w3329 & w3335;
	assign w3345 = w3344 & w3313;
	assign w3342 = w3341 ? w3293 : s420;
	assign w3341 = w3340 & w3313;
	assign w3340 = w3318 & w3335;
	assign w3552 = {63'b000000000000000000000000000000000000000000000000000000000000000, w23};
	assign w3338 = w3337 ? w3293 : s419;
	assign w3337 = w3336 & w3313;
	assign w3392 = w3391 & w3313;
	assign w3336 = w3302 & w3335;
	assign w4428 = w3831 & w4375;
	assign w3335 = w3334 & w3309;
	assign w3332 = w3331 ? w3293 : s418;
	assign w3331 = w3330 & w3313;
	assign w3330 = w3329 & w3310;
	assign w3329 = w3317 & w3323;
	assign w3327 = w3326 ? w3293 : s417;
	assign w3346 = w3345 ? w3293 : s421;
	assign w3326 = w3325 & w3313;
	assign w3325 = w3324 & w3310;
	assign w3324 = w3299 & w3323;
	assign w3323 = w3300 == w23;
	assign w4417 = w4416 & w3756;
	assign w3321 = w3320 ? w3293 : s416;
	assign w3320 = w3319 & w3313;
	assign w3319 = w3318 & w3310;
	assign w3317 = w3298 == w23;
	assign w3315 = w3314 ? w3293 : s415;
	assign w3314 = w3311 & w3313;
	assign w3313 = i12 ? w3312 : w47;
	assign w3312 = w299 ? w23 : w47;
	assign w3309 = w3306 & w3308;
	assign w3308 = w3307 == w47;
	assign w3306 = w3305 == w47;
	assign w3305 = w3297[3:3];
	assign w4797 = w4796 ? w3726 : s1986;
	assign w3303 = w3297[2:2];
	assign w3302 = w3299 & w3301;
	assign w3300 = w3297[1:1];
	assign w3299 = w3298 == w47;
	assign w3298 = w3297[0:0];
	assign w3297 = i12 ? w3296 : i40;
	assign w3296 = w299 ? w398 : i41;
	assign w3750 = w3731[7:7];
	assign w3417 = w3416 & w3313;
	assign w3286 = {15'b000000000000000, w1105};
	assign w3283 = s404 + w3282;
	assign w3282 = {15'b000000000000000, w1101};
	assign w4386 = w4385 ? w3726 : s1788;
	assign w3280 = i13 ? s305 : w117;
	assign w3278 = i12 ? w3277 : s297;
	assign w3277 = i13 ? w3276 : w47;
	assign w4762 = w3841 & w4701;
	assign w3276 = w982 ? w3275 : s297;
	assign w3273 = w3187 ? s297 : w3272;
	assign w4800 = w4799 & w3756;
	assign w3272 = w3184 ? w47 : s297;
	assign w3271 = w3177 ? w3270 : s297;
	assign w3270 = w294 ? w47 : s297;
	assign w3268 = w1453 ? w23 : w47;
	assign w3266 = w3265 ? w688 : w3262;
	assign w3265 = w3263 | w3264;
	assign w3263 = ~i13;
	assign w3256 = w3255 ? w3253 : w3252;
	assign w3254 = {3'b000, w23};
	assign w3253 = w2746 ? s180 : w23;
	assign w3252 = w3251 ? w3249 : s180;
	assign w4682 = w4681 & w3756;
	assign w3251 = s2760 == w3250;
	assign w4562 = w3836 & w4505;
	assign w3773 = w3772 ? w3726 : s1496;
	assign w3248 = w913 ? w47 : s180;
	assign w3246 = i13 ? w3245 : w47;
	assign w3245 = s2995 ? w3244 : w47;
	assign w3486 = w3459 ? s471 : s470;
	assign w3244 = w3243 ? s152 : w3241;
	assign w3242 = {2'b00, w44};
	assign w3241 = w3240 ? s152 : w3239;
	assign w3239 = w3238 ? w23 : s152;
	assign w3238 = ~w3237;
	assign w3237 = |s2997;
	assign w3231 = i12 ? w3230 : s121;
	assign w4708 = w4707 ? w3726 : s1945;
	assign w3230 = i13 ? w3229 : w47;
	assign w3229 = w982 ? w3228 : w23;
	assign w3228 = w3227 ? w23 : s121;
	assign w3226 = {1'b0, w44};
	assign w3224 = i13 ? w3223 : w117;
	assign w3222 = w2642 & s2632;
	assign w3220 = i13 ? w2532 : w696;
	assign w4094 = w4093 & w3756;
	assign w3215 = i13 ? w3214 : w47;
	assign w3213 = w3212 ? w3210 : w3207;
	assign w3212 = |w3211;
	assign w3210 = s55 ? w3209 : w23;
	assign w3485 = w3459 ? s469 : s468;
	assign w3207 = w3181 ? w3206 : s55;
	assign w4305 = w4304 & w3756;
	assign w3206 = w294 ? w47 : s55;
	assign w3637 = {w3636, w3635};
	assign w3201 = w902 ? w1028 : s31;
	assign w3199 = i12 ? w3198 : s22;
	assign w3197 = w982 ? w3196 : s22;
	assign w3195 = ~w3194;
	assign w4964 = s3000[31:31];
	assign w3559 = i13 ? w3558 : w1042;
	assign w3194 = |s2760;
	assign w3318 = w3317 & w3301;
	assign w3193 = s55 ? w3188 : w34;
	assign w3191 = s2760 == w3190;
	assign w3190 = {2'b00, w34};
	assign w3189 = s55 ? w3188 : w3183;
	assign w3187 = s55 & w3186;
	assign w4624 = w3831 & w4571;
	assign w3186 = ~w294;
	assign w3488 = w3459 ? s473 : s472;
	assign w3185 = w3184 ? w688 : s22;
	assign w3184 = s55 & w294;
	assign w3183 = {w47, w2763};
	assign w4943 = w3243 ? w4942 : w4940;
	assign w3182 = w3181 ? w3175 : s22;
	assign w3181 = |w3180;
	assign w3180 = {w3179, w3177};
	assign w3179 = s2760 == w3178;
	assign w3178 = {1'b0, w74};
	assign w3176 = {1'b0, w88};
	assign w3940 = w3793 & w3915;
	assign w3175 = w294 ? w688 : s22;
	assign w3172 = i12 ? w3171 : s18;
	assign w3169 = w3168 ? w3167 : w3152;
	assign w3168 = w398[4:4];
	assign w3167 = w3151 ? w3166 : w3159;
	assign w3164 = w3134 ? s475 : s474;
	assign w3163 = w3134 ? s473 : s472;
	assign w3162 = w3137 ? w3161 : w3160;
	assign w4109 = w3841 & w4048;
	assign w3361 = w3360 ? w3293 : s438;
	assign w3161 = w3134 ? s471 : s470;
	assign w3160 = w3134 ? s469 : s468;
	assign w3443 = w3302 & w3442;
	assign w3159 = w3142 ? w3158 : w3155;
	assign w3157 = w3134 ? s460 : s459;
	assign w3156 = w3134 ? s458 : s457;
	assign w3155 = w3137 ? w3154 : w3153;
	assign w3154 = w3134 ? s456 : s455;
	assign w3153 = w3134 ? s454 : s453;
	assign w3508 = w775 ? w791 : w3507;
	assign w3152 = w3151 ? w3150 : w3143;
	assign w3151 = w398[3:3];
	assign w3170 = |w398;
	assign w3149 = w3137 ? w3148 : w3147;
	assign w3148 = w3134 ? s444 : s443;
	assign w3147 = w3134 ? s442 : s441;
	assign w3146 = w3137 ? w3145 : w3144;
	assign w3145 = w3134 ? s440 : s439;
	assign w3144 = w3134 ? s438 : s437;
	assign w3143 = w3142 ? w3141 : w3138;
	assign w3138 = w3137 ? w3136 : w3135;
	assign w3137 = w398[1:1];
	assign w3451 = w3324 & w3442;
	assign w3135 = w3134 ? s416 : s415;
	assign w3134 = w398[0:0];
	assign w3132 = w629;
	assign w3131 = w655;
	assign w3130 = w668;
	assign w3781 = w3737 == w23;
	assign w3128 = w624;
	assign w3126 = w609;
	assign w3124 = w625;
	assign w3123 = w661;
	assign w3120 = w668;
	assign w3118 = w617;
	assign w3117 = w620;
	assign w3115 = w679;
	assign w3114 = w604;
	assign w4256 = w3776 & w4243;
	assign w3113 = w640;
	assign w4915 = w2746 ? w44 : w4914;
	assign w3112 = w574;
	assign w4940 = w3240 ? w4939 : s2997;
	assign w3110 = w580;
	assign w3109 = w631;
	assign w3108 = w634;
	assign w3105 = w654;
	assign w3103 = w651;
	assign w3223 = w2714 ? w3222 : w117;
	assign w3102 = w568;
	assign w3100 = w591;
	assign w3099 = w637;
	assign w4706 = w3762 & w4701;
	assign w3098 = i9;
	assign w3097 = w552;
	assign w4891 = i13 ? w4890 : w47;
	assign w3096 = w556;
	assign w3094 = i11[31:20];
	assign w3093 = w549;
	assign w3089 = w549;
	assign w4344 = w4343 & w3756;
	assign w3088 = w546;
	assign w3087 = w543;
	assign w3085 = s152;
	assign w3084 = s762;
	assign w3083 = s18;
	assign w3078 = w237;
	assign w3077 = w884;
	assign w3075 = s19;
	assign w3074 = s180;
	assign w3073 = s127;
	assign w3071 = i9;
	assign w3816 = w3815 & w3753;
	assign w3070 = w964;
	assign w3069 = s3011;
	assign w3067 = s2999;
	assign w4397 = w4396 & w3756;
	assign w3064 = w3063;
	assign w3063 = w963 ? w3062 : w3061;
	assign w3062 = s960[31:0];
	assign w3060 = w3059 ? s2971 : w3057;
	assign w3059 = |w3058;
	assign w3058 = {w217, w214};
	assign w3057 = w3056 ? s3011 : w3054;
	assign w3056 = |w3055;
	assign w3717 = ~w1441;
	assign w3618 = i13 ? w3617 : w3584;
	assign w3055 = {w211, w208};
	assign w3054 = w3053 ? s2991 : w3051;
	assign w3052 = {w205, w202};
	assign w3719 = w3717 + w3718;
	assign w3051 = w3050 ? s3047 : w3044;
	assign w3127 = w676;
	assign w3050 = |w3049;
	assign w3046 = s3045 & w1067;
	assign w3044 = w3043 ? s3040 : w3037;
	assign w4519 = w4518 & w3756;
	assign w3042 = {w196, w190};
	assign w4903 = w294 ? w42 : w88;
	assign w3039 = s3038 & w1067;
	assign w3036 = |w3035;
	assign w3711 = w1310 ? w3710 : w3707;
	assign w3035 = {w859, w3034};
	assign w4390 = w4389 ? w3726 : s1789;
	assign w3493 = w760[4:4];
	assign w3032 = {w851, w3031};
	assign w3028 = {w172, w169};
	assign w3027 = w3026 ? s3001 : w3024;
	assign w3984 = w3983 ? w3726 : s1591;
	assign w3026 = |w3025;
	assign w3025 = {w165, w162};
	assign w3092 = w556;
	assign w3022 = {w158, w156};
	assign w3020 = s2991;
	assign w3018 = w949;
	assign w3681 = s1294[34:1];
	assign w3014 = w951;
	assign w3012 = s960;
	assign w3010 = i9;
	assign w3009 = w944;
	assign w3008 = i13;
	assign w3007 = s18;
	assign w3004 = w944;
	assign w3003 = i13;
	assign w3002 = s18;
	assign w2998 = i9;
	assign w2992 = s18;
	assign w4982 = i13 ? w4981 : w117;
	assign w2988 = i13;
	assign w2987 = s18;
	assign w2986 = w945;
	assign w2985 = i9;
	assign w2984 = w944;
	assign w2979 = w944;
	assign w2978 = i13;
	assign w2976 = w951;
	assign w2975 = i9;
	assign w2974 = w944;
	assign w2973 = i13;
	assign w2972 = s18;
	assign w2970 = i9;
	assign w2968 = i13;
	assign w2966 = i9;
	assign w2964 = i13;
	assign w2963 = s18;
	assign w2962 = w760;
	assign w4264 = w3788 & w4243;
	assign w2961 = w376;
	assign w2960 = w397;
	assign w3188 = w3187 ? s22 : w3185;
	assign w2959 = s305;
	assign w2958 = w2957;
	assign w2956 = |w2955;
	assign w2952 = 12'b000000000000;
	assign w2951 = w368 ? w2950 : w2920;
	assign w2950 = {w2949, w2948};
	assign w2949 = s305[31:31];
	assign w2947 = s305[31:31];
	assign w2943 = s305[31:31];
	assign w2939 = s305[31:31];
	assign w2938 = {w2937, w2936};
	assign w2936 = {w2935, w2934};
	assign w3438 = w3329 & w3425;
	assign w2934 = {w2933, w2932};
	assign w2933 = s305[31:31];
	assign w2932 = {w2931, w2930};
	assign w2931 = s305[31:31];
	assign w2930 = {w2929, w2928};
	assign w2928 = {w2927, w2926};
	assign w2927 = s305[31:31];
	assign w2925 = s305[19:12];
	assign w2923 = s305[20:20];
	assign w2921 = s305[30:21];
	assign w3794 = w3793 & w3753;
	assign w2920 = w365 ? w2919 : w2918;
	assign w3535 = w3251 ? w3534 : s900;
	assign w2919 = w319 ? w2812 : w2767;
	assign w4120 = w4119 ? w3726 : s1657;
	assign w2917 = w359 ? w2916 : w2767;
	assign w3753 = w3747 & w3752;
	assign w2916 = {w2915, w2914};
	assign w2915 = s305[31:31];
	assign w2914 = {w2913, w2912};
	assign w2913 = s305[31:31];
	assign w2912 = {w2911, w2910};
	assign w2911 = s305[31:31];
	assign w2909 = s305[31:31];
	assign w4002 = w3788 & w3981;
	assign w2907 = s305[31:31];
	assign w4945 = i13 ? w4944 : w367;
	assign w3822 = w3821 & w3756;
	assign w2906 = {w2905, w2904};
	assign w4324 = w4323 & w3756;
	assign w2905 = s305[31:31];
	assign w2904 = {w2903, w2902};
	assign w2901 = s305[31:31];
	assign w2895 = s305[31:31];
	assign w2892 = {w2891, w2890};
	assign w2891 = s305[31:31];
	assign w2890 = {w2889, w2888};
	assign w2889 = s305[31:31];
	assign w4340 = w4339 & w3756;
	assign w3558 = w902 ? w3557 : s1011;
	assign w2888 = {w2887, w2886};
	assign w2886 = {w2885, w2884};
	assign w2885 = s305[31:31];
	assign w2884 = {w2883, w2882};
	assign w3080 = w944;
	assign w2883 = s305[31:31];
	assign w2882 = {w2881, w2880};
	assign w2878 = {w2877, w2876};
	assign w2875 = s305[7:7];
	assign w2873 = s305[30:25];
	assign w3525 = w3265 ? w688 : w3524;
	assign w2869 = w352 ? w2812 : w2767;
	assign w2868 = w348 ? w2867 : w2823;
	assign w2867 = w344 ? w2866 : w2767;
	assign w2863 = s305[31:31];
	assign w1273 = {w23, w1272};
	assign w3090 = w560;
	assign w222 = {w193, w221};
	assign w3171 = w3170 ? w3169 : w117;
	assign w2982 = s18;
	assign w1949 = w1494 ? s1948 : s1947;
	assign w1267 = w1130 ? w34 : w688;
	assign w1265 = i13;
	assign w1263 = w1237;
	assign w4872 = s2600 ? s2618 : w117;
	assign w4508 = w4507 ? w3726 : s1848;
	assign w3360 = w3359 & w3313;
	assign w1260 = w1259;
	assign w1259 = w1227[1:1];
	assign w2187 = i6;
	assign w1258 = w1257;
	assign w68 = |w67;
	assign w4493 = w3831 & w4440;
	assign w1213 = w1212 ? w1211 : w1206;
	assign w4511 = w4510 & w3756;
	assign w1205 = s1201 == w34;
	assign w976 = ~w975;
	assign w1253 = w1252;
	assign w518 = w516 & w517;
	assign w2587 = s31;
	assign w1980 = w1494 ? s1979 : s1978;
	assign w2216 = {w2215, w2214};
	assign w3690 = w3689 ? w3683 : i44;
	assign w595 = w594 & w558;
	assign w2690 = {6'b000000, w143};
	assign w1097 = i12;
	assign w4253 = w4252 & w3756;
	assign w3482 = w3459 ? s460 : s459;
	assign w1236 = 36'b000000000000000000000000000000000000;
	assign w4662 = w4661 & w3756;
	assign w1235 = s1234[36:1];
	assign w1228 = w1227;
	assign w569 = w563 | w568;
	assign w2896 = {w2895, w2894};
	assign w546 = i11[19:15];
	assign w1227 = w1220 ? w44 : w1226;
	assign w816 = s815;
	assign w1219 = |s1201;
	assign w818 = i12;
	assign w657 = i11[31:30];
	assign w353 = w352 ? w307 : w301;
	assign w1215 = s1201 == w1214;
	assign w1212 = s1201 == w32;
	assign w759 = w319 ? w367 : w301;
	assign w1210 = w1209 ? w23 : w47;
	assign w4219 = w3815 & w4178;
	assign w3141 = w3137 ? w3140 : w3139;
	assign w823 = w151;
	assign w3106 = w599;
	assign w1286 = i9;
	assign w873 = {w205, w871};
	assign w1202 = i13;
	assign w3748 = w3731[6:6];
	assign w1161 = s1160[34:1];
	assign w1194 = w1192 + w1193;
	assign w837 = {w832, w836};
	assign w3471 = w3462 ? w3470 : w3469;
	assign w1312 = w1289[0:0];
	assign w1192 = ~s1191;
	assign w3136 = w3134 ? s418 : s417;
	assign w1911 = w1525 ? w1910 : w1895;
	assign w3372 = w3302 & w3371;
	assign w3258 = i13 ? w3257 : w47;
	assign w2205 = i6[31:31];
	assign w4274 = w4273 ? w3726 : s1730;
	assign w1220 = ~w1219;
	assign w912 = s239 & w840;
	assign w1177 = w1176;
	assign w1176 = {w47, w1175};
	assign w4779 = w3776 & w4766;
	assign w203 = 10'b1100010011;
	assign w4540 = w4539 ? w3726 : s1863;
	assign w727 = w348 ? w726 : w725;
	assign w1173 = w1172 ? w1171 : w1168;
	assign w4507 = w4506 & w3756;
	assign w1167 = s762[30:0];
	assign w1872 = w1494 ? s1871 : s1870;
	assign w4057 = w3770 & w4048;
	assign w1163 = w1153[2:2];
	assign w4881 = w4858 ? w117 : w4880;
	assign w4102 = w4101 & w3756;
	assign w1126 = w299;
	assign w2630 = s2606;
	assign w3072 = w956;
	assign w1162 = 34'b0000000000000000000000000000000000;
	assign w4750 = w3826 & w4701;
	assign w1422 = {w1421, w1420};
	assign w1152 = w1141 ? w88 : w1151;
	assign w1151 = w1138 ? w74 : w42;
	assign w2140 = w2013[29:20];
	assign w1144 = {w47, w1143};
	assign w391 = w348 ? w390 : w389;
	assign w949 = ($signed(s18) < $signed(w944));
	assign w1142 = w1141 ? w32 : w1139;
	assign w4124 = w4123 ? w3726 : s1659;
	assign w1693 = w1494 ? s1692 : s1691;
	assign w4639 = w4638 ? w3726 : s1912;
	assign w1139 = w1138 ? w1137 : w1133;
	assign w1137 = {w23, w1136};
	assign w1136 = w1135 ? w23 : w47;
	assign w2224 = {w2223, w2222};
	assign w2777 = s305[31:31];
	assign w4389 = w4388 & w3756;
	assign w955 = w857 ? w954 : w953;
	assign w496 = w488[95:64];
	assign w1123 = s762;
	assign w377 = s305[11:7];
	assign w4932 = s18 | w944;
	assign w3810 = w3761 & w3804;
	assign w996 = w84;
	assign w1121 = s18;
	assign w1120 = w299;
	assign w3414 = w3413 ? w3293 : s458;
	assign w466 = {s459, w465};
	assign w1107 = w770;
	assign w1105 = w1104 ? w23 : w47;
	assign w4548 = w4547 ? w3726 : s1866;
	assign w3607 = w3604[16:16];
	assign w2780 = {w2779, w2778};
	assign w744 = s305[24:20];
	assign w3903 = w3902 ? w3726 : s1550;
	assign w1104 = w1098 & w1103;
	assign w1102 = w1101;
	assign w486 = w47 ? w451 : w436;
	assign w1101 = w1100 ? w23 : w47;
	assign w4086 = w4085 & w3756;
	assign w3490 = w3462 ? w3489 : w3488;
	assign w1100 = w1098 & w1099;
	assign w1098 = w401 & w299;
	assign w301 = 5'b11111;
	assign w3576 = {4'b0000, w23};
	assign w1092 = w299;
	assign w1091 = i13;
	assign w921 = {w196, w920};
	assign w2715 = w2714;
	assign w1089 = w1088;
	assign w1048 = s19 == w1047;
	assign w326 = |w325;
	assign w2576 = w278 ? w2561 : w2575;
	assign w2965 = w944;
	assign w2446 = {w2445, w2444};
	assign w4193 = w4192 ? w3726 : s1692;
	assign w2752 = w2748 == w2751;
	assign w1084 = w142 ? w1015 : w1083;
	assign w4546 = w3815 & w4505;
	assign w1079 = w151;
	assign w51 = s49 == w50;
	assign w2813 = w309 ? w2812 : w2767;
	assign w2696 = s19;
	assign w1078 = w151;
	assign w1077 = s815;
	assign w1420 = {w1419, w1418};
	assign w2028 = w2013[23:20];
	assign w1075 = w47;
	assign w4920 = w3179 ? w4919 : w4917;
	assign w3378 = w3377 ? w3293 : s442;
	assign w2955 = {w372, w370};
	assign w30 = w29 ? w20 : i14;
	assign w4097 = w3826 & w4048;
	assign w1074 = s19;
	assign w3561 = {63'b000000000000000000000000000000000000000000000000000000000000000, w23};
	assign w537 = w535 & w536;
	assign w1073 = w902;
	assign w3622 = i13 ? w3621 : w3620;
	assign w1068 = s1066 & w1067;
	assign w4796 = w4795 & w3756;
	assign w2657 = w2649 == w2656;
	assign w1065 = w1064;
	assign w3600 = w3597[16:16];
	assign w2775 = s305[31:31];
	assign w2481 = i6[15:15];
	assign w1434 = {w1433, w1432};
	assign w1060 = s1007[63:32];
	assign w73 = s49 == w72;
	assign w3724 = w802 ? w2012 : i45;
	assign w1056 = 12'b110000000000;
	assign w2519 = i8;
	assign w2766 = w736;
	assign w1164 = w1163 ? w1162 : w1161;
	assign w4636 = w3847 & w4570;
	assign w3598 = s1160[17:1];
	assign w1526 = w1525 ? w1524 : w1509;
	assign w2515 = w972 ? w2514 : w2511;
	assign w1054 = w1053 ? w1050 : w1049;
	assign w3420 = w3329 & w3407;
	assign w685 = i12 | w684;
	assign w1436 = {w1435, w1434};
	assign w2758 = i13;
	assign w4518 = w3776 & w4505;
	assign w1051 = 12'b110010000001;
	assign w700 = {w696, w699};
	assign w1376 = w1297[33:33];
	assign w1049 = w1048 ? w1045 : w1041;
	assign w175 = {w165, w174};
	assign w3311 = w3302 & w3310;
	assign w1252 = {w47, w1251};
	assign w1047 = {20'b00000000000000000000, w1046};
	assign w1041 = w1040 ? w1037 : w1036;
	assign w467 = {s460, w466};
	assign w1040 = s19 == w1039;
	assign w4498 = w4497 & w3756;
	assign w2989 = w944;
	assign w1038 = 12'b110010000010;
	assign w1532 = w1494 ? s1531 : s1530;
	assign w1216 = w1215 ? w32 : w1213;
	assign w1037 = s1011[63:32];
	assign w1036 = w1035 ? w1032 : w117;
	assign w283 = w244 ? w47 : w23;
	assign w2424 = {w2423, w2422};
	assign w1027 = w1026 ? w1016 : w1024;
	assign w3140 = w3134 ? s422 : s421;
	assign w1024 = w134 ? w1023 : w1022;
	assign w718 = s305[14:12];
	assign w1231 = i9;
	assign w318 = |w308;
	assign w2145 = w2027;
	assign w1017 = w1016;
	assign w4142 = w3798 & w4113;
	assign w1013 = {29'b00000000000000000000000000000, w44};
	assign w2573 = w51 ? w2572 : w2566;
	assign w4677 = w3815 & w4636;
	assign w3949 = w3948 & w3756;
	assign w1122 = w376;
	assign w1002 = w45;
	assign w1001 = i3;
	assign w1000 = w61;
	assign w777 = ~i2;
	assign w3445 = w3444 ? w3293 : s472;
	assign w2099 = w2046;
	assign w998 = w69;
	assign w631 = w630 & w628;
	assign w632 = w629 | w631;
	assign w997 = i4;
	assign w413 = w408 & w412;
	assign w992 = i6;
	assign w3999 = w3998 & w3756;
	assign w1605 = w1508 ? w1604 : w1597;
	assign w3805 = w3736 & w3804;
	assign w986 = w115;
	assign w3765 = w3764 ? w3726 : s1491;
	assign w3660 = w3659 ? w3657 : w3652;
	assign w3121 = w671;
	assign w681 = ~w23;
	assign w985 = s984;
	assign w3133 = w563;
	assign w719 = {w718, w717};
	assign w4808 = w4807 & w3756;
	assign w2579 = w80 ? w2578 : w696;
	assign w4372 = w4371 & w3756;
	assign w981 = w29 ? w980 : i21;
	assign w980 = w979 ? w978 : w973;
	assign w3086 = w543;
	assign w2317 = {w2316, w2315};
	assign w4189 = w4188 ? w3726 : s1691;
	assign w2429 = i6[31:31];
	assign w3758 = w3757 ? w3726 : s1490;
	assign w211 = s127 == w210;
	assign w548 = w545 & w547;
	assign w2068 = w2013[6:0];
	assign w4958 = w3240 ? w4957 : w4956;
	assign w2247 = {w2245, w2246};
	assign w2456 = i6[15:15];
	assign w969 = w968 ? w47 : w23;
	assign w968 = w20[0:0];
	assign w4011 = w4010 & w3756;
	assign w3669 = i13 ? w3668 : w3613;
	assign w966 = w293;
	assign w2046 = w2013[14:12];
	assign w3013 = s2971;
	assign w2593 = s762;
	assign w384 = w337 ? w383 : w382;
	assign w4490 = w4489 & w3756;
	assign w958 = i9;
	assign w228 = {w211, w227};
	assign w2311 = {w2310, w2309};
	assign w953 = w854 ? w952 : w950;
	assign w4715 = w4714 & w3756;
	assign w56 = w54 & s55;
	assign w952 = ~w951;
	assign w4301 = w4300 & w3756;
	assign w951 = s18 == w944;
	assign w950 = w851 ? w949 : w948;
	assign w947 = w845 ? w946 : w47;
	assign w245 = w244 ? w23 : w47;
	assign w945 = s18 < w944;
	assign w1197 = w1196;
	assign w1366 = w1326 + w1365;
	assign w2025 = |w2018;
	assign w941 = {w214, w940};
	assign w2662 = w2649 == w2661;
	assign w2410 = {w2408, w2409};
	assign w280 = w76 ? w279 : w268;
	assign w930 = {w854, w929};
	assign w2495 = w254 ? w117 : w2494;
	assign w1185 = {w835, w826};
	assign w1238 = w1237 ? w1236 : w1235;
	assign w929 = {w851, w928};
	assign w928 = {w848, w845};
	assign w926 = |w925;
	assign w1296 = w1289[2:2];
	assign w760 = w365 ? w759 : w758;
	assign w920 = {w169, w919};
	assign w911 = w151 | w887;
	assign w2586 = i12;
	assign w2588 = w811;
	assign w1275 = w1274 ? w1273 : w1269;
	assign w2346 = i6[15:15];
	assign w66 = {w33, w65};
	assign w4216 = w4215 & w3756;
	assign w3377 = w3376 & w3313;
	assign w536 = |s404;
	assign w908 = s55;
	assign w2673 = w2672 ? w2669 : w2668;
	assign w904 = s180;
	assign w247 = w56 ? w245 : w47;
	assign w1554 = w1494 ? s1553 : s1552;
	assign w903 = w902;
	assign w895 = s19;
	assign w3684 = s1294[1:0];
	assign w570 = {2'b00, w23};
	assign w891 = w890;
	assign w1206 = w1205 ? w1204 : i23;
	assign w1319 = {{2{w1297[33:33]}}, w1297};
	assign w890 = ~w889;
	assign w639 = w625 & w601;
	assign w888 = w887;
	assign w1240 = w1174[31:16];
	assign w886 = &s885;
	assign w3636 = s1234[36:36];
	assign w2698 = s127;
	assign w3807 = w3806 & w3756;
	assign w2980 = i9;
	assign w1138 = s1127 == w32;
	assign w1214 = {1'b0, w23};
	assign w359 = w331 | w358;
	assign w3744 = w3743 == w47;
	assign w407 = ~w406;
	assign w4897 = i10[31:2];
	assign w884 = w883 ? s180 : w842;
	assign w4007 = w4006 & w3756;
	assign w1083 = w138 ? s19 : w117;
	assign w871 = {w202, w870};
	assign w2737 = w736;
	assign w870 = {w199, w869};
	assign w893 = s305;
	assign w2059 = {w2058, w2057};
	assign w3614 = w1174[31:16];
	assign w1045 = s1043[31:0];
	assign w867 = {w190, w866};
	assign w4828 = w4827 & w3756;
	assign w2877 = s305[31:31];
	assign w869 = {w196, w868};
	assign w866 = {w186, w865};
	assign w865 = {w183, w864};
	assign w861 = {w851, w860};
	assign w1854 = w1499 ? w1853 : w1850;
	assign w855 = 10'b1011100011;
	assign w1190 = w1189;
	assign w1225 = w1212 ? w74 : w42;
	assign w3594 = |w3593;
	assign w961 = s960[32:32];
	assign w972 = w737 == w971;
	assign w854 = s127 == w853;
	assign w4245 = w4244 & w3756;
	assign w853 = {4'b0000, w852};
	assign w171 = {2'b00, w170};
	assign w2651 = {7'b0000000, w2650};
	assign w849 = 10'b1001100011;
	assign w848 = s127 == w847;
	assign w847 = {2'b00, w846};
	assign w3893 = w3820 & w3848;
	assign w846 = 10'b1101100011;
	assign w1943 = w1558 ? w1942 : w1911;
	assign w4959 = s3000[31:4];
	assign w2127 = {w2126, w2125};
	assign w3869 = w3788 & w3848;
	assign w844 = {2'b00, w843};
	assign w4313 = w4312 ? w3726 : s1754;
	assign w1099 = w398 < w544;
	assign w1950 = w1499 ? w1949 : w1946;
	assign w2497 = i7;
	assign w3431 = w3430 & w3313;
	assign w835 = s127 == w834;
	assign w831 = {1'b0, w830};
	assign w830 = 11'b10110110011;
	assign w3729 = w802 ? w3728 : i47;
	assign w1014 = s31 + w1013;
	assign w829 = s127 == w828;
	assign w1025 = s127[6:0];
	assign w824 = 11'b10010110011;
	assign w198 = {3'b000, w197};
	assign w2922 = {w2921, w47};
	assign w822 = w237;
	assign w594 = w551 & w593;
	assign w2842 = {w2841, w2840};
	assign w2367 = i6[7:7];
	assign w3889 = w3815 & w3848;
	assign w3497 = i12 ? w3496 : s762;
	assign w821 = w255;
	assign w4884 = w2714 ? w2644 : w4883;
	assign w1257 = w1255 + w1256;
	assign w2881 = s305[31:31];
	assign w2256 = i6[23:23];
	assign w820 = w151;
	assign w263 = w73 ? w262 : w257;
	assign w2161 = w2012;
	assign w2248 = w974 == w34;
	assign w3478 = w3459 ? s454 : s453;
	assign w817 = s31;
	assign w814 = s813;
	assign w1112 = w760;
	assign w1132 = s1127 == w34;
	assign w812 = w811;
	assign w1953 = w1494 ? s1952 : s1951;
	assign w809 = ~w808;
	assign w2924 = {w2923, w2922};
	assign w807 = w804 & w806;
	assign w3752 = w3749 & w3751;
	assign w806 = ~w805;
	assign w2237 = i6[31:31];
	assign w4131 = w4130 & w3756;
	assign w3620 = 17'b00000000000000000;
	assign w805 = s792 == s797;
	assign w1809 = w1494 ? s1808 : s1807;
	assign w1247 = w1187[31:16];
	assign w1917 = w1494 ? s1916 : s1915;
	assign w37 = |w36;
	assign w3628 = w1261 ? w3627 : s1207;
	assign w796 = w794 + w795;
	assign w3709 = {w3708, w47};
	assign w1241 = {1'b0, w1240};
	assign w1165 = w1164;
	assign w795 = {7'b0000000, w23};
	assign w1297 = w1296 ? w1162 : w1295;
	assign w4538 = w3805 & w4505;
	assign w1072 = i9;
	assign w785 = w29 ? w47 : i19;
	assign w291 = w56 ? w283 : w290;
	assign w2910 = {w2909, w2908};
	assign w783 = w778 & w782;
	assign w1750 = w1558 ? w1749 : w1718;
	assign w781 = w780 == w678;
	assign w3198 = i13 ? w3197 : w688;
	assign w1279 = w1130 ? w23 : w47;
	assign w779 = 6'b000000;
	assign w2241 = {w2240, w2239};
	assign w774 = s772;
	assign w771 = w770;
	assign w1469 = s18;
	assign w770 = w234 ? s769 : i18;
	assign w767 = w397;
	assign w1646 = w1499 ? w1645 : w1642;
	assign w765 = s18;
	assign w763 = s762;
	assign w653 = w649 & w566;
	assign w2385 = i6[7:7];
	assign w957 = w956;
	assign w1262 = w1261;
	assign w758 = w362 ? w757 : w756;
	assign w1179 = {w47, w1178};
	assign w563 = w559 & w562;
	assign w2865 = s305[31:31];
	assign w1683 = w1494 ? s1682 : s1681;
	assign w3538 = w982 ? w3537 : s900;
	assign w946 = ~w945;
	assign w2397 = i6[7:7];
	assign w1145 = |s1127;
	assign w3806 = w3805 & w3753;
	assign w230 = {w217, w229};
	assign w757 = w359 ? w744 : w301;
	assign w2149 = w2095;
	assign w753 = w344 ? w744 : w301;
	assign w752 = w388 ? w367 : w751;
	assign w1211 = {w23, w1210};
	assign w3122 = w551;
	assign w321 = w311 == w143;
	assign w803 = ~w802;
	assign w381 = w319 ? w377 : w380;
	assign w1412 = w1297[33:33];
	assign w2691 = w2649 == w2690;
	assign w750 = w334 ? w744 : w301;
	assign w3890 = w3889 & w3756;
	assign w2554 = w266 ? w86 : w2553;
	assign w749 = w321 ? w748 : w746;
	assign w3104 = w596;
	assign w860 = {w848, w845};
	assign w1523 = w1499 ? w1522 : w1519;
	assign w939 = {w202, w938};
	assign w1339 = {w1337, w1336};
	assign w745 = w309 ? w744 : w301;
	assign w3139 = w3134 ? s420 : s419;
	assign w1157 = i9;
	assign w4304 = w3841 & w4243;
	assign w756 = w355 ? w755 : w754;
	assign w742 = w741;
	assign w739 = s121;
	assign w934 = {w158, w933};
	assign w1759 = w1494 ? s1758 : s1757;
	assign w737 = w736[8:7];
	assign w209 = 10'b1000010011;
	assign w1250 = {1'b0, w1249};
	assign w1860 = w1494 ? s1859 : s1858;
	assign w480 = {s473, w479};
	assign w2154 = w2013;
	assign w4901 = 4'b0100;
	assign w892 = i11;
	assign w1059 = w1058 ? w1055 : w1054;
	assign w736 = w375 ? w735 : w733;
	assign w251 = w25 ? w250 : i17;
	assign w1676 = w1494 ? s1675 : s1674;
	assign w2181 = w38;
	assign w1080 = s127;
	assign w3654 = s1234[18:1];
	assign w3101 = w676;
	assign w863 = {w857, w862};
	assign w4288 = w3820 & w4243;
	assign w2228 = {w2227, w2226};
	assign w1416 = {w1415, w1414};
	assign w728 = w352 ? w692 : w687;
	assign w726 = w344 ? w692 : w687;
	assign w2055 = w2054 ? w2020 : w2052;
	assign w723 = w722 ? w720 : w716;
	assign w596 = w595 & w562;
	assign w3037 = w3036 ? w117 : w3030;
	assign w964 = w963 ? w961 : w47;
	assign w720 = {w47, w719};
	assign w1015 = s31 + s19;
	assign w1125 = i13;
	assign w715 = s305[30:30];
	assign w4948 = {w47, w4947};
	assign w2123 = w2013[14:12];
	assign w3262 = {w3261, w234};
	assign w975 = |w974;
	assign w2507 = s762[7:0];
	assign w1992 = w1494 ? s1991 : s1990;
	assign w970 = s55 ? w969 : w23;
	assign w330 = w328 == w329;
	assign w1284 = w1283;
	assign w2552 = w264 ? w42 : w88;
	assign w4720 = w4719 ? w3726 : s1951;
	assign w1147 = w1146 ? w1144 : w1142;
	assign w710 = w334 ? w709 : w687;
	assign w3715 = i13 ? w3714 : w3620;
	assign w2431 = i6[31:31];
	assign w1149 = s1134;
	assign w2370 = {w2369, w2368};
	assign w706 = s305[25:25];
	assign w948 = w848 ? w945 : w947;
	assign w1239 = w1238;
	assign w1932 = w1494 ? s1931 : s1930;
	assign w2494 = w25 ? w2493 : i26;
	assign w1096 = w401;
	assign w3996 = w3995 ? w3726 : s1595;
	assign w764 = w376;
	assign w1649 = w1494 ? s1648 : s1647;
	assign w711 = w337 ? w710 : w702;
	assign w2294 = i6[23:23];
	assign w3107 = w586;
	assign w2658 = w2657 ? w2654 : w2653;
	assign w2590 = w255;
	assign w705 = {w704, w703};
	assign w2013 = w802 ? w2012 : w2010;
	assign w702 = w321 ? w701 : w694;
	assign w4418 = w4417 ? w3726 : s1803;
	assign w1733 = w1508 ? w1732 : w1725;
	assign w1103 = w398 >= w544;
	assign w910 = w294;
	assign w701 = w319 ? w700 : w695;
	assign w699 = {w698, w697};
	assign w4329 = w4328 ? w3726 : s1761;
	assign w550 = w549 < w544;
	assign w693 = w309 ? w692 : w687;
	assign w1131 = w1130 ? w34 : w688;
	assign w2730 = s18;
	assign w691 = {w690, w689};
	assign w2208 = {w2207, w2206};
	assign w2589 = w770;
	assign w690 = s305[14:12];
	assign w1418 = {w1417, w1416};
	assign w2425 = i6[31:31];
	assign w4416 = w3815 & w4375;
	assign w2693 = w2692[7:7];
	assign w2266 = i6[23:23];
	assign w1665 = w1494 ? s1664 : s1663;
	assign w680 = w677 | w679;
	assign w679 = w560 == w678;
	assign w1108 = i9;
	assign w4315 = w3762 & w4310;
	assign w624 = w621 | w623;
	assign w4449 = w3770 & w4440;
	assign w2453 = w2452 ? w2451 : i32;
	assign w672 = w671 & w663;
	assign w670 = w659 & w545;
	assign w350 = s305[14:13];
	assign w4393 = w4392 & w3756;
	assign w4095 = w4094 ? w3726 : s1644;
	assign w3274 = s55 ? w3273 : w2763;
	assign w3214 = w982 ? w3213 : s55;
	assign w669 = w656 | w668;
	assign w991 = i7;
	assign w4534 = w3798 & w4505;
	assign w2926 = {w2925, w2924};
	assign w2085 = {w2084, w2083};
	assign w3150 = w3142 ? w3149 : w3146;
	assign w664 = w661 & w663;
	assign w3974 = w3973 ? w3726 : s1585;
	assign w663 = ~w662;
	assign w660 = w659 & w547;
	assign w1200 = w1163;
	assign w2050 = w2049 ? w2042 : w2013;
	assign w2093 = w2092;
	assign w656 = w624 | w655;
	assign w194 = 9'b110010011;
	assign w2591 = i13;
	assign w655 = w652 | w654;
	assign w1424 = {w1423, w1422};
	assign w3410 = w3409 ? w3293 : s457;
	assign w2395 = i6[7:7];
	assign w3453 = w3452 ? w3293 : s474;
	assign w2711 = w2710;
	assign w1154 = w1153;
	assign w1251 = w1248 + w1250;
	assign w647 = w646 & w628;
	assign w4164 = w4163 ? w3726 : s1678;
	assign w889 = &s127;
	assign w324 = s305[31:31];
	assign w322 = w321 ? w320 : w315;
	assign w2582 = w244 ? s49 : w2581;
	assign w320 = w319 ? w307 : w317;
	assign w2121 = w2013[6:0];
	assign w1050 = s1043[63:32];
	assign w1124 = w760;
	assign w3708 = w1174[15:0];
	assign w365 = w311 == w132;
	assign w583 = w552 == w582;
	assign w356 = w355 ? w353 : w349;
	assign w666 = w560 == w665;
	assign w1481 = |w1480;
	assign w3356 = w3355 & w3313;
	assign w1918 = w1499 ? w1917 : w1914;
	assign w2653 = w2652 ? w2648 : w2647;
	assign w4861 = w4846 ? w23 : w47;
	assign w1119 = w397;
	assign w313 = {2'b00, w312};
	assign w1128 = i13;
	assign w2714 = w2692[6:6];
	assign w909 = s239;
	assign w310 = w309 ? w307 : w301;
	assign w169 = s127 == w168;
	assign w3307 = w3297[4:4];
	assign w676 = w675 & w577;
	assign w530 = w528 & w529;
	assign w614 = w613 & w562;
	assign w309 = |w308;
	assign w2072 = {w2027, w2071};
	assign w1245 = {w47, w1244};
	assign w922 = {w199, w921};
	assign w826 = s127 == w825;
	assign w1274 = s1264 == w32;
	assign w2222 = {w2221, w2220};
	assign w603 = w602 & w558;
	assign w304 = s302 & w303;
	assign w4634 = w4633 ? w3726 : s1907;
	assign w1608 = w1494 ? s1607 : s1606;
	assign w303 = 32'b00000000000000000000000001111111;
	assign w651 = w650 & w628;
	assign w2058 = w2013[14:12];
	assign w2434 = {w2433, w2432};
	assign w819 = s118;
	assign w1968 = w1494 ? s1967 : s1966;
	assign w2555 = w90 ? w2554 : w2551;
	assign w311 = s305[6:0];
	assign w3158 = w3137 ? w3157 : w3156;
	assign w277 = ~i8;
	assign w94 = |w93;
	assign w709 = {w708, w707};
	assign w543 = i11[24:20];
	assign w786 = w37 ? w23 : w785;
	assign w3743 = w3731[4:4];
	assign w832 = s127 == w831;
	assign w79 = w78 ? w23 : w47;
	assign w1229 = w1130;
	assign w973 = w972 ? w970 : w23;
	assign w285 = w272 ? w23 : w47;
	assign w1965 = w1499 ? w1964 : w1961;
	assign w678 = 7'b1111111;
	assign w3691 = s1294[34:18];
	assign w3125 = w643;
	assign w842 = w178 ? s152 : w47;
	assign w221 = {w190, w220};
	assign w588 = w552 == w44;
	assign w278 = i4 & w277;
	assign w516 = w514 & w515;
	assign w897 = s896;
	assign w2872 = {w2871, w47};
	assign w172 = s127 == w171;
	assign w372 = w311 == w371;
	assign w712 = s305[6:0];
	assign w358 = ~w357;
	assign w2261 = {w2260, w2259};
	assign w988 = i8;
	assign w1187 = w1186 ? w1184 : s18;
	assign w1924 = w1494 ? s1923 : s1922;
	assign w2095 = w2013[31:20];
	assign w2703 = w2642;
	assign w266 = i8 & w260;
	assign w2825 = s305[31:25];
	assign w3621 = w1196 ? w1189 : s1191;
	assign w244 = i3 & i7;
	assign w117 = 32'b00000000000000000000000000000000;
	assign w857 = s127 == w856;
	assign w265 = w264 ? w47 : w23;
	assign w510 = w488[223:192];
	assign w1387 = {w1385, w1384};
	assign w1071 = w956;
	assign w4180 = w4179 & w3756;
	assign w3249 = w2754 ? w47 : w3248;
	assign w246 = w51 ? w245 : w243;
	assign w2420 = {w2419, w2418};
	assign w182 = {6'b000000, w181};
	assign w300 = w125 & w299;
	assign w615 = w610 | w614;
	assign w2344 = i6[15:15];
	assign w424 = {s416, s415};
	assign w2114 = w805;
	assign w1662 = w1499 ? w1661 : w1658;
	assign w3447 = w3318 & w3442;
	assign w463 = {s456, w462};
	assign w1053 = s19 == w1052;
	assign w293 = i13 ? w292 : w47;
	assign w264 = i8 & i5;
	assign w192 = {3'b000, w191};
	assign w1198 = w1153[0:0];
	assign w4990 = i13 ? w949 : w47;
	assign w623 = w622 & w562;
	assign w1249 = w1187[15:0];
	assign w258 = i4 & i5;
	assign w255 = w254 ? w47 : w251;
	assign w1093 = i13;
	assign w254 = |w253;
	assign w2441 = i6[31:31];
	assign w2462 = {w2461, w2460};
	assign w2634 = w2633 ? w47 : w23;
	assign w243 = w100 ? w242 : w47;
	assign w4302 = w4301 ? w3726 : s1744;
	assign w3656 = w3653[17:17];
	assign w1905 = w1494 ? s1904 : s1903;
	assign w956 = w859 ? w951 : w955;
	assign w3902 = w3901 & w3756;
	assign w883 = |w882;
	assign w646 = w645 & w558;
	assign w199 = s127 == w198;
	assign w919 = {w162, w918};
	assign w3359 = w3318 & w3354;
	assign w242 = i7 ? w23 : w47;
	assign w248 = w59 ? w247 : w246;
	assign w308 = s305[14:12];
	assign w1111 = w398;
	assign w2196 = {w2195, w2194};
	assign w267 = w266 ? w23 : w265;
	assign w619 = w578 & w612;
	assign w227 = {w208, w226};
	assign w299 = w296 & w298;
	assign w1465 = w840;
	assign w571 = w552 == w570;
	assign w1826 = w1494 ? s1825 : s1824;
	assign w3720 = w1473 ? w3719 : w1441;
	assign w2837 = s305[31:31];
	assign w226 = {w205, w225};
	assign w4791 = w3793 & w4766;
	assign w2185 = i5;
	assign w477 = {s470, w476};
	assign w1326 = {w1325, w117};
	assign w2309 = {w2308, w2307};
	assign w999 = w38;
	assign w485 = w484[31:0];
	assign w223 = {w196, w222};
	assign w3918 = w3917 ? w3726 : s1560;
	assign w2723 = s118;
	assign w2981 = w949;
	assign w538 = w537 & w401;
	assign w1109 = w760;
	assign w218 = 12'b100000110011;
	assign w509 = w506 & w508;
	assign w270 = w269 & i5;
	assign w3815 = w3769 & w3804;
	assign w1623 = s1492[5:5];
	assign w216 = {2'b00, w215};
	assign w272 = w269 & w260;
	assign w462 = {s455, w461};
	assign w1438 = {w1437, w1436};
	assign w214 = s127 == w213;
	assign w4610 = w4609 ? w3726 : s1897;
	assign w2315 = {w2314, w2313};
	assign w3467 = w760[2:2];
	assign w1581 = w1499 ? w1580 : w1577;
	assign w3549 = w2710 ? s18 : w3548;
	assign w1369 = w1297[33:33];
	assign w2078 = w2013[6:0];
	assign w1061 = 12'b110010000000;
	assign w4038 = w3836 & w3981;
	assign w307 = s305[19:15];
	assign w3393 = w3392 ? w3293 : s453;
	assign w141 = {7'b0000000, w140};
	assign w4019 = w4018 & w3756;
	assign w1226 = w1215 ? w88 : w1225;
	assign w599 = w598 & w562;
	assign w27 = ~w26;
	assign w4074 = w4073 & w3756;
	assign w704 = s305[14:12];
	assign w3528 = w2638 ? w23 : w3527;
	assign w207 = {2'b00, w206};
	assign w3749 = w3748 == w47;
	assign w2641 = w47;
	assign w3803 = w3739 == w23;
	assign w1116 = s18;
	assign w4433 = w4432 & w3756;
	assign w206 = 10'b1000110011;
	assign w4865 = s2611 ? w47 : s2612;
	assign w2321 = {w2320, w2319};
	assign w253 = {w35, w252};
	assign w2056 = w2013[6:0];
	assign w2473 = i6[15:15];
	assign w2568 = i3 & w2567;
	assign w3367 = w3329 & w3354;
	assign w696 = 4'b0000;
	assign w20 = s18 + s19;
	assign w987 = s109;
	assign w3871 = w3870 ? w3726 : s1535;
	assign w426 = {s417, w424};
	assign w2467 = i6[15:15];
	assign w3496 = w3495 ? w3494 : w117;
	assign w579 = w578 & w558;
	assign w4361 = w4360 ? w3726 : s1776;
	assign w2115 = w800;
	assign w4503 = w4502 ? w3726 : s1843;
	assign w3569 = {31'b0000000000000000000000000000000, w23};
	assign w347 = {1'b0, w346};
	assign w3204 = i13 ? w2584 : w696;
	assign w197 = 9'b100010011;
	assign w262 = w261 ? w23 : w259;
	assign w925 = {w217, w924};
	assign w1555 = w1499 ? w1554 : w1551;
	assign w386 = {w370, w385};
	assign w2749 = {1'b0, w346};
	assign w138 = s127 == w137;
	assign w4825 = w4824 ? w3726 : s2000;
	assign w90 = s49 == w89;
	assign w4771 = w3762 & w4766;
	assign w74 = 3'b101;
	assign w2414 = w2413 ? w2411 : w117;
	assign w3982 = w3742 & w3981;
	assign w312 = 5'b11000;
	assign w414 = ~w413;
	assign w1857 = w1494 ? s1856 : s1855;
	assign w882 = {w219, w880};
	assign w833 = 11'b10100110011;
	assign w1411 = {w1409, w1408};
	assign w661 = w660 & w550;
	assign w82 = w56 ? w47 : w81;
	assign w1868 = w1494 ? s1867 : s1866;
	assign w4970 = i13 ? w4969 : w117;
	assign w76 = s49 == w75;
	assign w506 = w502 & w505;
	assign w213 = {2'b00, w212};
	assign w2817 = {w2815, w2816};
	assign w513 = s422 == s460;
	assign w493 = w491 == w492;
	assign w1086 = |w1085;
	assign w1752 = s1492[6:6];
	assign w1875 = w1494 ? s1874 : s1873;
	assign w1182 = w1180 + w1181;
	assign w69 = w68 ? w42 : i16;
	assign w158 = s127 == w157;
	assign w284 = w51 ? w283 : w282;
	assign w688 = 2'b00;
	assign w1507 = w1499 ? w1506 : w1503;
	assign w177 = {w172, w176};
	assign w2439 = i6[31:31];
	assign w559 = w555 & w558;
	assign w4138 = w3793 & w4113;
	assign w2835 = s305[31:31];
	assign w931 = {w857, w930};
	assign w3624 = i13 ? w1221 : w688;
	assign w1133 = w1132 ? w1131 : i22;
	assign w3068 = s3006;
	assign w649 = w625 & w593;
	assign w2776 = {w2775, w2774};
	assign w4200 = w4199 & w3756;
	assign w366 = w365 ? w364 : w363;
	assign w2879 = s305[31:31];
	assign w249 = i13 ? w248 : w47;
	assign w3465 = w3459 ? s422 : s421;
	assign w261 = i4 & w260;
	assign w44 = 3'b100;
	assign w4675 = w4674 ? w3726 : s1928;
	assign w71 = 3'b111;
	assign w733 = w365 ? w732 : w731;
	assign w1118 = w770;
	assign w937 = {w190, w936};
	assign w1787 = w1494 ? s1786 : s1785;
	assign w4764 = w4763 ? w3726 : s1970;
	assign w1005 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
	assign w3662 = 19'b0000000000000000000;
	assign w181 = 6'b110011;
	assign w3546 = i13 ? w3545 : w3542;
	assign w983 = w982;
	assign w2134 = {w2133, w2132};
	assign w668 = w667 & w577;
	assign w2263 = {w2262, w2261};
	assign w643 = w642 & w628;
	assign w2789 = s305[31:31];
	assign w1524 = w1508 ? w1523 : w1516;
	assign w155 = {1'b0, w154};
	assign w378 = w309 ? w377 : w301;
	assign w4555 = w4554 & w3756;
	assign w2541 = w786;
	assign w609 = w608 & w562;
	assign w78 = |w77;
	assign w4847 = w4846 ? w117 : w4845;
	assign w290 = w80 ? w289 : w47;
	assign w36 = {w35, w33};
	assign w1290 = w1289;
	assign w2583 = w56 ? w2582 : w2579;
	assign w3029 = |w3028;
	assign w271 = w270 ? w47 : w23;
	assign w160 = 8'b10010011;
	assign w1886 = w1494 ? s1885 : s1884;
	assign w3202 = i13 ? w3201 : w117;
	assign w2652 = w2649 == w2651;
	assign w3243 = s2997 >= w3242;
	assign w478 = {s471, w477};
	assign w4473 = w3805 & w4440;
	assign w151 = w150 ? w23 : w47;
	assign w191 = 9'b100110011;
	assign w3866 = w3865 & w3756;
	assign w174 = {w162, w173};
	assign w1218 = {w47, w1217};
	assign w3499 = i13 ? w3063 : w117;
	assign w2953 = s305[31:12];
	assign w183 = s127 == w182;
	assign w582 = {1'b0, w34};
	assign w810 = w803 & w809;
	assign w4951 = {w696, w4950};
	assign w29 = |w28;
	assign w880 = {w217, w878};
	assign w388 = |w387;
	assign w1620 = w1508 ? w1619 : w1612;
	assign w137 = {6'b000000, w136};
	assign w3579 = ~i13;
	assign w273 = w272 ? w23 : w271;
	assign w487 = w47 ? w482 : w467;
	assign w2272 = i6[23:23];
	assign w535 = s404 == s409;
	assign w1209 = s1207 == w1208;
	assign w4050 = w4049 & w3756;
	assign w185 = {7'b0000000, w184};
	assign w648 = w644 | w647;
	assign w2592 = s18;
	assign w286 = w275 ? w23 : w285;
	assign w163 = 8'b10110011;
	assign w445 = {s438, s437};
	assign w789 = ~w788;
	assign w994 = i5;
	assign w4252 = w3770 & w4243;
	assign w42 = 3'b000;
	assign w4987 = i13 ? w945 : w47;
	assign w2941 = s305[31:31];
	assign w776 = ~w775;
	assign w54 = w53 | w25;
	assign w4010 = w3798 & w3981;
	assign w238 = w151 | w237;
	assign w3424 = w3352 & w3388;
	assign w1815 = w1525 ? w1814 : w1799;
	assign w3412 = w3318 & w3407;
	assign w1087 = w1086 ? w1014 : w1084;
	assign w907 = s180;
	assign w4375 = w3847 & w4309;
	assign w1199 = w1198;
	assign w327 = ~w326;
	assign w355 = w311 == w354;
	assign w3116 = w623;
	assign w586 = w585 & w562;
	assign w84 = i13 ? w83 : w47;
	assign w3119 = w614;
	assign w2550 = w261 ? w86 : w2549;
	assign w936 = {w172, w935};
	assign w2413 = ~w2412;
	assign w2639 = w2638;
	assign w979 = w737 == w32;
	assign w52 = w51 ? w23 : w47;
	assign w282 = w100 ? w281 : w280;
	assign w4969 = s2995 ? w4968 : s18;
	assign w4568 = w4567 ? w3726 : s1874;
	assign w1499 = s1492[1:1];
	assign w219 = s127 == w218;
	assign w1148 = w1147;
	assign w836 = {w829, w826};
	assign w590 = w589 & w558;
	assign w2942 = {w2941, w2940};
	assign w1006 = s1004 & w1005;
	assign w26 = |s22;
	assign w3755 = w802 ? w23 : w47;
	assign w1697 = w1494 ? s1696 : s1695;
	assign w977 = w976 ? w23 : w47;
	assign w3240 = |s2997;
	assign w1242 = w1174[15:0];
	assign w176 = {w169, w175};
	assign w354 = {5'b00000, w34};
	assign w1794 = w1494 ? s1793 : s1792;
	assign w641 = w638 | w640;
	assign w4281 = w4280 & w3756;
	assign w149 = {w145, w148};
	assign w2683 = w2682 ? w2679 : w2678;
	assign w794 = {1'b0, s792};
	assign w93 = {w76, w92};
	assign w4430 = w4429 ? w3726 : s1808;
	assign w566 = w556 == w565;
	assign w2801 = s305[31:31];
	assign w4978 = s2995 ? w4977 : s18;
	assign w1169 = ~s762;
	assign w802 = w790 & w801;
	assign w4694 = w4693 & w3756;
	assign w645 = w625 & w571;
	assign w2113 = w2009;
	assign w1174 = w826 ? w1173 : s762;
	assign w593 = w552 == w74;
	assign w2659 = 9'b001000000;
	assign w233 = |w232;
	assign w1237 = w1227[2:2];
	assign w1276 = {1'b0, w23};
	assign w1146 = ~w1145;
	assign w722 = w342 != w721;
	assign w3586 = s1160[34:1];
	assign w150 = |w149;
	assign w104 = w59 ? w57 : w103;
	assign w2572 = {w688, w2571};
	assign w95 = w94 ? w23 : w47;
	assign w989 = s107;
	assign w725 = w340 ? w724 : w711;
	assign w45 = w37 ? w44 : w43;
	assign w1340 = w1328[33:33];
	assign w2283 = {w2282, w2281};
	assign w4098 = w4097 & w3756;
	assign w1035 = s19 == w1034;
	assign w791 = 7'b0000000;
	assign w340 = w311 == w339;
	assign w677 = w669 | w676;
	assign w2042 = {w2033, w2041};
	assign w465 = {s458, w464};
	assign w240 = w238 | s239;
	assign w1890 = w1494 ? s1889 : s1888;
	assign w1181 = {31'b0000000000000000000000000000000, w23};
	assign w281 = i7 ? w47 : w23;
	assign w574 = w573 & w562;
	assign w993 = w105;
	assign w489 = w488[31:0];
	assign w1716 = w1499 ? w1715 : w1712;
	assign w4528 = w4527 ? w3726 : s1856;
	assign w878 = {w214, w876};
	assign w2745 = w736 == w2744;
	assign w1717 = w1508 ? w1716 : w1709;
	assign w2637 = |i10;
	assign w2654 = 9'b010000000;
	assign w2768 = s305[31:20];
	assign w698 = s305[20:20];
	assign w1117 = s762;
	assign w342 = s305[13:12];
	assign w298 = s180 | s297;
	assign w189 = {3'b000, w188};
	assign w344 = w332 & w343;
	assign w630 = w625 & w577;
	assign w24 = {1'b0, w23};
	assign w4512 = w4511 ? w3726 : s1849;
	assign w1224 = i9;
	assign w59 = ~w58;
	assign w2067 = w2066 ? w2063 : w2050;
	assign w2623 = i9;
	assign w990 = s22;
	assign w1168 = {w47, w1167};
	assign w514 = w512 & w513;
	assign w3264 = ~s180;
	assign w3091 = i11;
	assign w47 = 1'b0;
	assign w2672 = w2649 == w2671;
	assign w4727 = w4726 & w3756;
	assign w287 = w278 ? w23 : w286;
	assign w2903 = s305[31:31];
	assign w2621 = s2606;
	assign w202 = s127 == w201;
	assign w3349 = w3348 & w3313;
	assign w1639 = w1508 ? w1638 : w1631;
	assign w3216 = i12 ? w3215 : s55;
	assign w621 = w618 | w620;
	assign w2969 = w944;
	assign w2091 = w2043;
	assign w775 = ~i12;
	assign w373 = {w370, w368};
	assign w1999 = w1494 ? s1998 : s1997;
	assign w2259 = {w2258, w2257};
	assign w4965 = {w4964, w4963};
	assign w3936 = w3788 & w3915;
	assign w751 = w337 ? w750 : w749;
	assign w236 = &s235;
	assign w1437 = w1297[33:33];
	assign w96 = w59 ? w82 : w95;
	assign w858 = {5'b00000, w361};
	assign w721 = {1'b0, w23};
	assign w633 = w625 & w583;
	assign w1055 = s1007[31:0];
	assign w611 = {6'b000000, w23};
	assign w2253 = {w2252, w2251};
	assign w102 = |w101;
	assign w4310 = w3747 & w4309;
	assign w81 = w80 ? w23 : w47;
	assign w1483 = w1482;
	assign w1156 = i13;
	assign w852 = 8'b11100011;
	assign w2017 = w2014;
	assign w370 = w311 == w369;
	assign w1052 = {20'b00000000000000000000, w1051};
	assign w205 = s127 == w204;
	assign w1088 = w145 ? w1064 : w1087;
	assign w577 = w552 == w576;
	assign w606 = w552 == w71;
	assign w3732 = w3731[0:0];
	assign w1450 = ~w1237;
	assign w35 = s22 == w34;
	assign w4008 = w4007 ? w3726 : s1601;
	assign w58 = |s49;
	assign w279 = w278 ? w23 : w276;
	assign w2280 = i6[23:23];
	assign w131 = s127 == w130;
	assign w2773 = s305[31:31];
	assign w1668 = w1494 ? s1667 : s1666;
	assign w1942 = w1525 ? w1941 : w1926;
	assign w4894 = i13 ? w4893 : w117;
	assign w4257 = w4256 & w3756;
	assign w2839 = s305[31:31];
	assign w4738 = w3810 & w4701;
	assign w1184 = w1183 ? w1182 : w1179;
	assign w707 = {w706, w705};
	assign w184 = 5'b10011;
	assign w1030 = w1014;
	assign w2538 = w293;
	assign w552 = i11[14:12];
	assign w1031 = w1015;
	assign w4212 = w4211 & w3756;
	assign w2016 = w775;
	assign w97 = i13 ? w96 : w47;
	assign w3647 = s1234[18:1];
	assign w1141 = s1127 == w1140;
	assign w112 = |w111;
	assign w557 = |w556;
	assign w503 = w484[159:128];
	assign w1336 = {w1334, w1333};
	assign w292 = w59 ? w291 : w284;
	assign w1183 = s18[31:31];
	assign w1522 = w1494 ? s1521 : s1520;
	assign w2469 = i6[15:15];
	assign w87 = s49 == w86;
	assign w674 = w560 == w673;
	assign w367 = 5'b00000;
	assign w2996 = s2995;
	assign w1208 = 5'b10001;
	assign w2977 = s18;
	assign w613 = w555 & w612;
	assign w288 = w274 & w277;
	assign w4702 = w3742 & w4701;
	assign w4266 = w4265 ? w3726 : s1727;
	assign w1153 = w1146 ? w44 : w1152;
	assign w1150 = i9;
	assign w115 = i13 ? w114 : w47;
	assign w1417 = w1297[33:33];
	assign w4711 = w4710 & w3756;
	assign w839 = |w838;
	assign w99 = {2'b00, w34};
	assign w4090 = w4089 & w3756;
	assign w3384 = w3329 & w3371;
	assign w113 = w112 ? w23 : w47;
	assign w2339 = {w2338, w2337};
	assign w2372 = {w2371, w2370};
	assign w4494 = w4493 & w3756;
	assign w317 = w316 ? w307 : w301;
	assign w940 = {w208, w939};
	assign w259 = w258 ? w47 : w23;
	assign w2491 = w2490 ? w2489 : w2453;
	assign w1289 = w1282 ? w44 : w1288;
	assign w408 = w401 & w407;
	assign w2173 = w2043;
	assign w3808 = w3807 ? w3726 : s1510;
	assign w208 = s127 == w207;
	assign w4835 = i13 ? w4834 : w117;
	assign w3304 = w3303 == w47;
	assign w162 = s127 == w161;
	assign w1223 = s1207;
	assign w4550 = w3820 & w4505;
	assign w2533 = w2532;
	assign w4957 = s3000[31:1];
	assign w3399 = w3324 & w3390;
	assign w604 = w603 & w562;
	assign w2347 = {w2346, w2345};
	assign w133 = {5'b00000, w132};
	assign w2201 = i6[31:31];
	assign w341 = w340 ? w307 : w338;
	assign w260 = ~i5;
	assign w1221 = w1220 ? w1218 : w1216;
	assign w4544 = w4543 ? w3726 : s1864;
	assign w1621 = w1525 ? w1620 : w1605;
	assign w4954 = i13 ? w4953 : w117;
	assign w2479 = i6[15:15];
	assign w1189 = {w47, w1188};
	assign w105 = i13 ? w104 : w47;
	assign w2290 = i6[23:23];
	assign w580 = w579 & w562;
	assign w605 = w600 | w604;
	assign w2527 = 4'b1100;
	assign w1343 = w1328[33:33];
	assign w923 = {w205, w922};
	assign w111 = {w76, w90};
	assign w4469 = w3798 & w4440;
	assign w490 = w485 == w489;
	assign w335 = w334 ? w307 : w301;
	assign w4642 = w4641 & w3756;
	assign w4489 = w3826 & w4440;
	assign w1170 = {31'b0000000000000000000000000000000, w23};
	assign w447 = {s440, w446};
	assign w3177 = s2760 == w3176;
	assign w1638 = w1499 ? w1637 : w1634;
	assign w3520 = w47 ? s31 : s815;
	assign w2595 = w737;
	assign w887 = w884 & w886;
	assign w1441 = w1366 + w1440;
	assign w1178 = s18[30:0];
	assign w2856 = {w2855, w2854};
	assign w100 = s49 == w99;
	assign w2722 = w2721;
	assign w1268 = s1264 == w34;
	assign w2516 = w979 ? s762 : w2515;
	assign w3208 = w3184 ? w47 : w23;
	assign w499 = w484[127:96];
	assign w876 = {w211, w875};
	assign w274 = ~i4;
	assign w515 = s437 == s468;
	assign w545 = w543 < w544;
	assign w1486 = w1174;
	assign w125 = i0 & i12;
	assign w129 = 7'b1101111;
	assign w1311 = w1310;
	assign w132 = 7'b1100111;
	assign w4156 = w4155 ? w3726 : s1674;
	assign w1172 = s762[31:31];
	assign w2064 = {5'b00000, w34};
	assign w86 = 4'b1000;
	assign w50 = {2'b00, w32};
	assign w1313 = w1312;
	assign w3566 = w3565 ? w3562 : s1043;
	assign w140 = 5'b10111;
	assign w83 = w59 ? w82 : w79;
	assign w1280 = {w47, w1279};
	assign w3043 = |w3042;
	assign w2871 = s305[11:8];
	assign w2543 = s55;
	assign w3795 = w3794 & w3756;
	assign w393 = w355 ? w392 : w391;
	assign w1346 = w1328[33:33];
	assign w1244 = w1241 + w1243;
	assign w3920 = w3762 & w3915;
	assign w2614 = w2613;
	assign w2104 = w2087;
	assign w1480 = {w835, w1479};
	assign w215 = 10'b1110010011;
	assign w428 = {s418, w426};
	assign w3582 = w3581 ? w367 : w3578;
	assign w2990 = i9;
	assign w2302 = w974 == w32;
	assign w3492 = w3476 ? w3491 : w3484;
	assign w334 = w327 | w333;
	assign w766 = w299;
	assign w193 = s127 == w192;
	assign w2874 = {w2873, w2872};
	assign w1988 = w1499 ? w1987 : w1984;
	assign w1195 = w1194;
	assign w4869 = s2601 ? w47 : w2613;
	assign w2704 = s2632;
	assign w38 = w37 ? s31 : w30;
	assign w2004 = w1508 ? w2003 : w1996;
	assign w314 = w311 == w313;
	assign w4196 = w4195 & w3756;
	assign w1544 = w1494 ? s1543 : s1542;
	assign w1566 = w1499 ? w1565 : w1562;
	assign w210 = {2'b00, w209};
	assign w1435 = w1297[33:33];
	assign w2066 = w2065 & w2048;
	assign w1370 = {w1369, w1368};
	assign w157 = 12'b101010110011;
	assign w905 = s297;
	assign w636 = w625 & w588;
	assign w4816 = w4815 & w3756;
	assign w89 = {1'b0, w88};
	assign w2578 = w288 ? w2577 : w2576;
	assign w4906 = w3184 ? w696 : s2760;
	assign w3234 = i12 ? w3233 : w47;
	assign w165 = s127 == w164;
	assign w1799 = w1508 ? w1798 : w1791;
	assign w2558 = w272 ? w86 : w2557;
	assign w170 = 10'b1010110011;
	assign w561 = {1'b0, w181};
	assign w4053 = w3762 & w4048;
	assign w1539 = w1494 ? s1538 : s1537;
	assign w694 = w314 ? w693 : w687;
	assign w2605 = s2604 & w1067;
	assign w4703 = w4702 & w3756;
	assign w2733 = w47;
	assign w3081 = w770;
	assign w379 = w314 ? w378 : w301;
	assign w4481 = w3815 & w4440;
	assign w788 = ~w787;
	assign w2525 = w2413 ? w2524 : w696;
	assign w4653 = w3783 & w4636;
	assign w2567 = ~i7;
	assign w91 = {w73, w87};
	assign w4935 = w3265 ? w47 : s180;
	assign w808 = w807 & w789;
	assign w635 = w632 | w634;
	assign w3553 = s1007 + w3552;
	assign w713 = s305[14:12];
	assign w2361 = i6[7:7];
	assign w88 = 3'b110;
	assign w2994 = w944;
	assign w754 = w348 ? w753 : w752;
	assign w436 = {s422, w434};
	assign w178 = |w177;
	assign w33 = s22 == w32;
	assign w954 = ~w949;
	assign w57 = w56 ? w23 : w47;
	assign w154 = 11'b11010010011;
	assign w2098 = w2092;
	assign w3648 = {w3646, w3647};
	assign w1217 = w1130 ? w23 : w47;
	assign w2081 = {w2080, w2079};
	assign w3275 = w3191 ? w3274 : w3271;
	assign w612 = w556 == w611;
	assign w3870 = w3869 & w3756;
	assign w901 = w899 & s900;
	assign w1415 = w1297[33:33];
	assign w2218 = {w2217, w2216};
	assign w2751 = {5'b00000, w34};
	assign w1094 = i0;
	assign w1405 = {w1403, w1402};
	assign w3425 = w3304 & w3424;
	assign w828 = {1'b0, w827};
	assign w708 = s305[30:30];
	assign w782 = ~w781;
	assign w167 = 10'b1010010011;
	assign w186 = s127 == w185;
	assign w584 = w551 & w583;
	assign w1135 = s1134 == w544;
	assign w1603 = w1494 ? s1602 : s1601;
	assign w329 = {6'b000000, w23};
	assign w234 = w233 ? s180 : w179;
	assign w576 = {1'b0, w32};
	assign w332 = ~w331;
	assign w333 = w330 & w332;
	assign w387 = {w372, w386};
	assign w92 = {w90, w91};
	assign w755 = w352 ? w367 : w301;
	assign w3019 = w952;
	assign w894 = i10;
	assign w2360 = i6[7:7];
	assign w337 = w311 == w336;
	assign w4485 = w3820 & w4440;
	assign w2451 = {w2449, w2450};
	assign w671 = w670 & w547;
	assign w4351 = w3815 & w4310;
	assign w1457 = w1242;
	assign w4425 = w4424 & w3756;
	assign w338 = w337 ? w335 : w322;
	assign w1180 = ~s18;
	assign w345 = w344 ? w307 : w301;
	assign w2694 = w2634 & w2693;
	assign w61 = i13 ? w60 : w47;
	assign w1081 = s31;
	assign w1910 = w1508 ? w1909 : w1902;
	assign w252 = {w33, w27};
	assign w658 = |w657;
	assign w348 = w311 == w347;
	assign w1813 = w1499 ? w1812 : w1809;
	assign w2544 = s19;
	assign w1631 = w1499 ? w1630 : w1627;
	assign w3391 = w3302 & w3390;
	assign w662 = |w546;
	assign w913 = w911 | w912;
	assign w3065 = s3001;
	assign w2033 = 2'b01;
	assign w382 = w321 ? w381 : w379;
	assign w357 = |w350;
	assign w1488 = w811;
	assign w488 = w23 ? w487 : w486;
	assign w3033 = {w854, w3032};
	assign w491 = w484[63:32];
	assign w360 = w359 ? w307 : w301;
	assign w3456 = w3455 & w3313;
	assign w497 = w495 == w496;
	assign w2377 = i6[7:7];
	assign w734 = s305[6:0];
	assign w144 = {5'b00000, w143};
	assign w1451 = w1449 & w1450;
	assign w1454 = w1453;
	assign w3095 = w3094;
	assign w927 = w926 ? s19 : i20;
	assign w361 = 7'b1100011;
	assign w364 = w319 ? w307 : w301;
	assign w4426 = w4425 ? w3726 : s1807;
	assign w2097 = w2012;
	assign w1106 = w1105;
	assign w2324 = i6[15:15];
	assign w1033 = 12'b110000000010;
	assign w2898 = {w2897, w2896};
	assign w173 = {w158, w156};
	assign w368 = w311 == w129;
	assign w3440 = w3439 ? w3293 : s471;
	assign w1690 = w1494 ? s1689 : s1688;
	assign w1130 = s180 & w840;
	assign w2142 = w2013[29:25];
	assign w2482 = {w2481, w2480};
	assign w450 = {s443, w449};
	assign w942 = {w219, w941};
	assign w1292 = i13;
	assign w1893 = w1494 ? s1892 : s1891;
	assign w269 = i4 & i8;
	assign w375 = |w374;
	assign w995 = w97;
	assign w965 = w964;
	assign w3973 = w3972 & w3756;
	assign w3863 = w3862 ? w3726 : s1531;
	assign w3702 = w3699[16:16];
	assign w692 = {w688, w691};
	assign w1082 = w770;
	assign w380 = w316 ? w377 : w301;
	assign w1026 = w1025 == w361;
	assign w2450 = i6[31:16];
	assign w2740 = w902;
	assign w328 = s305[31:25];
	assign w4093 = w3820 & w4048;
	assign w3030 = w3029 ? s2999 : w3027;
	assign w1841 = w1494 ? s1840 : s1839;
	assign w389 = w388 ? w377 : w384;
	assign w1277 = s1264 == w1276;
	assign w4803 = w3810 & w4766;
	assign w2375 = i6[7:7];
	assign w3580 = s1134 == w544;
	assign w682 = w680 | w681;
	assign w294 = ~w293;
	assign w392 = w352 ? w377 : w301;
	assign w4849 = w4848 ? w4847 : s2606;
	assign w146 = {w134, w131};
	assign w899 = ~s898;
	assign w2401 = i6[7:7];
	assign w617 = w616 & w562;
	assign w3676 = s1270 == w544;
	assign w578 = w551 & w577;
	assign w4646 = w4645 & w3756;
	assign w638 = w635 | w637;
	assign w1333 = {w1331, w1330};
	assign w2929 = s305[31:31];
	assign w526 = w524 & w525;
	assign w2946 = {w2945, w2944};
	assign w1547 = w1494 ? s1546 : s1545;
	assign w394 = w359 ? w367 : w301;
	assign w346 = 6'b100011;
	assign w2726 = s813;
	assign w4294 = w4293 ? w3726 : s1741;
	assign w352 = w344 | w351;
	assign w3076 = w887;
	assign w397 = w365 ? w396 : w395;
	assign w4028 = w4027 ? w3726 : s1610;
	assign w53 = s22[1:1];
	assign w501 = w499 == w500;
	assign w1196 = w1153[1:1];
	assign w608 = w607 & w558;
	assign w2900 = {w2899, w2898};
	assign w732 = w319 ? w692 : w687;
	assign w2153 = w2088;
	assign w982 = w37 ? w23 : w981;
	assign w2275 = {w2274, w2273};
	assign w400 = w300 & w399;
	assign w1440 = {w1439, w1438};
	assign w406 = |s404;
	assign w1419 = w1297[33:33];
	assign w67 = {w35, w66};
	assign w383 = w334 ? w377 : w301;
	assign w411 = |s409;
	assign w840 = w839 ? w23 : w47;
	assign w1300 = {w47, w1299};
	assign w1515 = w1494 ? s1514 : s1513;
	assign w363 = w362 ? w360 : w356;
	assign w2048 = w2046 == w2047;
	assign w735 = {w367, w734};
	assign w412 = ~w411;
	assign w597 = w592 | w596;
	assign w3796 = w3795 ? w3726 : s1504;
	assign w2948 = {w2947, w2946};
	assign w190 = s127 == w189;
	assign w924 = {w211, w923};
	assign w1394 = w1297[33:33];
	assign w565 = {1'b0, w564};
	assign w4440 = w3914 & w4309;
	assign w430 = {s419, w428};
	assign w2918 = w362 ? w2917 : w2870;
	assign w1022 = w131 ? w1015 : w1021;
	assign w1003 = w38;
	assign w4497 = w3836 & w4440;
	assign w2069 = {w2055, w2068};
	assign w654 = w653 & w628;
	assign w1358 = w1328[33:33];
	assign w1278 = w1277 ? w32 : w1275;
	assign w492 = w488[63:32];
	assign w1034 = {20'b00000000000000000000, w1033};
	assign w1658 = w1494 ? s1657 : s1656;
	assign w1797 = w1494 ? s1796 : s1795;
	assign w432 = {s420, w430};
	assign w4420 = w3820 & w4375;
	assign w323 = s305[29:25];
	assign w4878 = {31'b0000000000000000000000000000000, w23};
	assign w3061 = w219 ? s3006 : w3060;
	assign w1887 = w1499 ? w1886 : w1883;
	assign w446 = {s439, w445};
	assign w452 = w47 ? w451 : w436;
	assign w4348 = w4347 & w3756;
	assign w554 = ~w553;
	assign w4363 = w3831 & w4310;
	assign w448 = {s441, w447};
	assign w4227 = w3826 & w4178;
	assign w2023 = w2013[18:15];
	assign w3257 = w982 ? w3256 : s180;
	assign w2815 = 20'b00000000000000000000;
	assign w3005 = i9;
	assign w2880 = {w2879, w2878};
	assign w1140 = {1'b0, w23};
	assign w75 = {1'b0, w74};
	assign w1042 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	assign w1021 = w1020 ? s815 : w1014;
	assign w2133 = w2013[29:25];
	assign w1476 = s1467[31:0];
	assign w3396 = w3395 & w3313;
	assign w449 = {s442, w448};
	assign w461 = {s454, s453};
	assign w747 = w316 ? w367 : w301;
	assign w906 = s180;
	assign w2688 = w2687 ? w2684 : w2683;
	assign w268 = w90 ? w267 : w263;
	assign w484 = w47 ? w483 : w452;
	assign w667 = w664 & w666;
	assign w2638 = w2637 ? w23 : w47;
	assign w4604 = w3805 & w4571;
	assign w494 = w490 & w493;
	assign w938 = {w193, w937};
	assign w834 = {1'b0, w833};
	assign w495 = w484[95:64];
	assign w601 = w552 == w88;
	assign w3721 = w1453 ? w3720 : w1042;
	assign w2402 = {w2401, w2400};
	assign w1956 = w1494 ? s1955 : s1954;
	assign w498 = w494 & w497;
	assign w652 = w648 | w651;
	assign w500 = w488[127:96];
	assign w164 = {4'b0000, w163};
	assign w390 = w344 ? w367 : w301;
	assign w1443 = w1440;
	assign w2087 = w2043 == w2086;
	assign w3688 = {w3687, w3685};
	assign w2243 = 24'b000000000000000000000000;
	assign w505 = w503 == w504;
	assign w628 = w560 == w627;
	assign w914 = w913;
	assign w23 = 1'b1;
	assign w602 = w551 & w601;
	assign w2565 = {w688, w2564};
	assign w2090 = s305;
	assign w508 = w507 == s458;
	assign w3474 = w3462 ? w3473 : w3472;
	assign w547 = w546 < w544;
	assign w220 = {w186, w183};
	assign w1751 = w1623 ? w1750 : w1687;
	assign w2041 = {w2039, w2038};
	assign w2260 = i6[23:23];
	assign w511 = s421 == w510;
	assign w512 = w509 & w511;
	assign w517 = s438 == s469;
	assign w1023 = s18 + s19;
	assign w1085 = {w134, w131};
	assign w2211 = i6[31:31];
	assign w520 = w518 & w519;
	assign w2386 = {w2385, w2384};
	assign w3933 = w3932 & w3756;
	assign w1782 = w1499 ? w1781 : w1778;
	assign w1261 = w1227[0:0];
	assign w521 = s440 == s471;
	assign w522 = w520 & w521;
	assign w2899 = s305[31:31];
	assign w902 = w901 ? w23 : w47;
	assign w3848 = w3847 & w3752;
	assign w3023 = |w3022;
	assign w1246 = w1245;
	assign w790 = w783 & w789;
	assign w1402 = {w1400, w1399};
	assign w528 = w526 & w527;
	assign w4357 = w4356 ? w3726 : s1773;
	assign w1186 = |w1185;
	assign w524 = w522 & w523;
	assign w1484 = w1187;
	assign w525 = s442 == s473;
	assign w527 = s443 == s474;
	assign w2112 = w802;
	assign w371 = {1'b0, w136};
	assign w385 = {w368, w340};
	assign w841 = w840;
	assign w531 = w414 | w530;
	assign w4744 = w4743 ? w3726 : s1962;
	assign w2144 = w2055;
	assign w1039 = {20'b00000000000000000000, w1038};
	assign w746 = w314 ? w745 : w301;
	assign w3839 = w3838 ? w3726 : s1520;
	assign w532 = ~w23;
	assign w591 = w590 & w562;
	assign w1357 = {w1355, w1354};
	assign w3785 = w3784 & w3756;
	assign w2859 = s305[31:31];
	assign w1028 = w47 ? s813 : w1027;
	assign w533 = w531 | w532;
	assign w3066 = s3000;
	assign w3034 = {w857, w3033};
	assign w1018 = 10'b1110011000;
	assign w864 = {w859, w863};
	assign w4981 = s18 - w944;
	assign w2459 = i6[15:15];
	assign w369 = {2'b00, w140};
	assign w541 = ~w540;
	assign w401 = s123 | w400;
	assign w2551 = w73 ? w2550 : w2547;
	assign w544 = 5'b10000;
	assign w697 = s305[6:0];
	assign w2129 = w2085;
	assign w549 = i11[11:7];
	assign w212 = 10'b1110110011;
	assign w3629 = s1207 == w1208;
	assign w551 = w548 & w550;
	assign w916 = s127;
	assign w4030 = w3826 & w3981;
	assign w761 = w760;
	assign w2022 = w2013;
	assign w555 = w551 & w554;
	assign w1677 = w1499 ? w1676 : w1673;
	assign w556 = i11[31:25];
	assign w3079 = w234;
	assign w560 = i11[6:0];
	assign w4491 = w4490 ? w3726 : s1839;
	assign w616 = w572 & w612;
	assign w3017 = w945;
	assign w567 = w555 & w566;
	assign w2276 = i6[23:23];
	assign w1171 = w1169 + w1170;
	assign w4272 = w3798 & w4243;
	assign w2314 = i6[15:15];
	assign w589 = w551 & w588;
	assign w1255 = ~s1254;
	assign w250 = w249 ? w23 : w47;
	assign w295 = w255 & w294;
	assign w932 = {w859, w931};
	assign w2782 = {w2781, w2780};
	assign w856 = {2'b00, w855};
	assign w572 = w551 & w571;
	assign w2111 = w2012;
	assign w3602 = w3589 == w32;
	assign w573 = w572 & w558;
	assign w114 = w59 ? w82 : w113;
	assign w575 = w569 | w574;
	assign w275 = w274 & i8;
	assign w581 = w575 | w580;
	assign w2465 = i6[15:15];
	assign w542 = w23 & w541;
	assign w1193 = {16'b0000000000000000, w23};
	assign w1654 = w1508 ? w1653 : w1646;
	assign w3737 = w3731[2:2];
	assign w587 = w581 | w586;
	assign w675 = w672 & w674;
	assign w399 = |w398;
	assign w598 = w594 & w566;
	assign w4114 = w3742 & w4113;
	assign w610 = w605 | w609;
	assign w729 = w355 ? w728 : w727;
	assign w974 = w20[1:0];
	assign w618 = w615 | w617;
	assign w620 = w619 & w562;
	assign w665 = {5'b00000, w34};
	assign w4244 = w3742 & w4243;
	assign w625 = w547 & w550;
	assign w2650 = 6'b110001;
	assign w2192 = i6[31:31];
	assign w336 = {1'b0, w181};
	assign w2862 = {w2861, w2860};
	assign w629 = w626 & w628;
	assign w4075 = w4074 ? w3726 : s1635;
	assign w130 = {5'b00000, w129};
	assign w1281 = |s1264;
	assign w2902 = {w2901, w2900};
	assign w257 = w87 ? w256 : w47;
	assign w2524 = w2522 << w2523;
	assign w963 = |w962;
	assign w4820 = w4819 & w3756;
	assign w2944 = {w2943, w2942};
	assign w343 = w342 != w34;
	assign w3442 = w3334 & w3424;
	assign w2034 = w2013[14:0];
	assign w592 = w587 | w591;
	assign w1375 = {w1373, w1372};
	assign w4815 = w3826 & w4766;
	assign w3862 = w3861 & w3756;
	assign w868 = {w193, w867};
	assign w634 = w633 & w628;
	assign w351 = w350 == w32;
	assign w237 = w234 & w236;
	assign w935 = {w165, w934};
	assign w2937 = s305[31:31];
	assign w1360 = {w1358, w1357};
	assign w147 = {w138, w146};
	assign w562 = w560 == w561;
	assign w4758 = w3836 & w4701;
	assign w640 = w639 & w628;
	assign w650 = w649 & w558;
	assign w1879 = w1558 ? w1878 : w1847;
	assign w2045 = w2043 == w2044;
	assign w743 = i13;
	assign w2509 = s762[7:0];
	assign w4404 = w3798 & w4375;
	assign w1282 = ~w1281;
	assign w2197 = i6[31:31];
	assign w2675 = 10'b1100110001;
	assign w1283 = w1282 ? w1280 : w1278;
	assign w4162 = w3826 & w4113;
	assign w644 = w641 | w643;
	assign w2217 = i6[31:31];
	assign w403 = 16'b0000000000000000;
	assign w1285 = s1270;
	assign w1110 = w398;
	assign w1287 = w1274 ? w74 : w42;
	assign w825 = {1'b0, w824};
	assign w1288 = w1277 ? w88 : w1287;
	assign w3502 = w982 ? w3501 : s772;
	assign w1291 = w1130;
	assign w1293 = i9;
	assign w2138 = w2087;
	assign w1298 = w1297;
	assign w196 = s127 == w195;
	assign w1557 = w1525 ? w1556 : w1541;
	assign w2834 = {w2833, w2832};
	assign w1299 = w1174[15:0];
	assign w1301 = w1300;
	assign w1302 = w1187[15:0];
	assign w3540 = i12 ? w3539 : s900;
	assign w1622 = w1558 ? w1621 : w1590;
	assign w2252 = i6[23:23];
	assign w1303 = {w47, w1302};
	assign w4691 = w4690 ? w3726 : s1935;
	assign w1304 = w1303;
	assign w1306 = ~s1305;
	assign w1307 = {16'b0000000000000000, w23};
	assign w1019 = {2'b00, w1018};
	assign w1455 = w1249;
	assign w3885 = w3810 & w3848;
	assign w2354 = i6[15:8];
	assign w1308 = w1306 + w1307;
	assign w1314 = w1296;
	assign w1316 = w1130;
	assign w1317 = w1252;
	assign w3111 = w647;
	assign w1320 = -w1319;
	assign w4823 = w3836 & w4766;
	assign w1321 = w1320;
	assign w1322 = {{2{w1164[33:33]}}, w1164};
	assign w4323 = w3776 & w4310;
	assign w2743 = 8'b11110011;
	assign w637 = w636 & w628;
	assign w1325 = w1164[31:0];
	assign w1328 = w1327 + w1320;
	assign w2368 = {w2367, w2366};
	assign w1331 = w1328[33:33];
	assign w4450 = w4449 & w3756;
	assign w2163 = w2076;
	assign w4571 = w3747 & w4570;
	assign w1095 = w537;
	assign w1512 = w1494 ? s1511 : s1510;
	assign w2049 = w2045 & w2048;
	assign w1342 = {w1340, w1339};
	assign w1345 = {w1343, w1342};
	assign w4844 = {31'b0000000000000000000000000000000, w23};
	assign w1348 = {w1346, w1345};
	assign w2026 = ~w2025;
	assign w1349 = w1328[33:33];
	assign w627 = {2'b00, w184};
	assign w1354 = {w1352, w1351};
	assign w3591 = |w3589;
	assign w1661 = w1494 ? s1660 : s1659;
	assign w1363 = {w1361, w1360};
	assign w4651 = w4650 ? w3726 : s1916;
	assign w1365 = {w1364, w1363};
	assign w1367 = w1297[33:33];
	assign w1368 = {w1367, w1297};
	assign w1371 = w1297[33:33];
	assign w3516 = s18 + s19;
	assign w2077 = w2076 ? w2074 : w2067;
	assign w1372 = {w1371, w1370};
	assign w943 = |w942;
	assign w1373 = w1297[33:33];
	assign w3364 = w3363 & w3313;
	assign w1378 = {w1376, w1375};
	assign w217 = s127 == w216;
	assign w1379 = w1297[33:33];
	assign w224 = {w199, w223};
	assign w2848 = {w2847, w2846};
	assign w4944 = s2995 ? w4943 : w4937;
	assign w3408 = w3302 & w3407;
	assign w1381 = {w1379, w1378};
	assign w1482 = w1481 ? w1478 : w1477;
	assign w1382 = w1297[33:33];
	assign w3608 = {w3607, w3606};
	assign w142 = s127 == w141;
	assign w2356 = {1'b0, w23};
	assign w1384 = {w1382, w1381};
	assign w2150 = w2020;
	assign w2732 = i13;
	assign w77 = {w76, w73};
	assign w1385 = w1297[33:33];
	assign w1894 = w1499 ? w1893 : w1890;
	assign w1390 = {w1388, w1387};
	assign w1391 = w1297[33:33];
	assign w2857 = s305[31:31];
	assign w1393 = {w1391, w1390};
	assign w2044 = {1'b0, w346};
	assign w1396 = {w1394, w1393};
	assign w1397 = w1297[33:33];
	assign w2870 = w355 ? w2869 : w2868;
	assign w395 = w362 ? w394 : w393;
	assign w1399 = {w1397, w1396};
	assign w3630 = w3579 | w3629;
	assign w1032 = s1011[31:0];
	assign w1400 = w1297[33:33];
	assign w1406 = w1297[33:33];
	assign w4685 = w3826 & w4636;
	assign w3233 = w299 ? i0 : s123;
	assign w1718 = w1525 ? w1717 : w1702;
	assign w2633 = |s2632;
	assign w1408 = {w1406, w1405};
	assign w4704 = w4703 ? w3726 : s1944;
	assign w464 = {s457, w463};
	assign w2610 = s2609;
	assign w1409 = w1297[33:33];
	assign w2183 = w84;
	assign w1421 = w1297[33:33];
	assign w1685 = w1508 ? w1684 : w1677;
	assign w1423 = w1297[33:33];
	assign w4609 = w4608 & w3756;
	assign w3823 = w3822 ? w3726 : s1514;
	assign w1462 = w1164;
	assign w1973 = w1508 ? w1972 : w1965;
	assign w2786 = {w2785, w2784};
	assign w3537 = w3255 ? w3536 : w3535;
	assign w626 = w625 & w554;
	assign w1426 = {w1425, w1424};
	assign w1427 = w1297[33:33];
	assign w1428 = {w1427, w1426};
	assign w4046 = w3748 == w23;
	assign w2051 = w2013[10:7];
	assign w1429 = w1297[33:33];
	assign w1432 = {w1431, w1430};
	assign w4960 = s3000[31:31];
	assign w2724 = s31;
	assign w2124 = {w2123, w2122};
	assign w4233 = w4232 ? w3726 : s1711;
	assign w1433 = w1297[33:33];
	assign w1439 = w1297[33:33];
	assign w3334 = w3303 == w23;
	assign w1442 = w1441;
	assign w2492 = w972 ? w2491 : w2414;
	assign w1444 = w1365;
	assign w1445 = w1326;
	assign w1446 = w1153;
	assign w553 = |w552;
	assign w1468 = i13;
	assign w4085 = w3810 & w4048;
	assign w2687 = w2649 == w2686;
	assign w862 = {w854, w861};
	assign w1447 = w1227;
	assign w714 = {w713, w712};
	assign w2531 = w979 ? w2530 : w2529;
	assign w1448 = w1289;
	assign w3981 = w3980 & w3752;
	assign w673 = {1'b0, w346};
	assign w1449 = ~w1163;
	assign w4014 = w3805 & w3981;
	assign w1452 = ~w1296;
	assign w3710 = {w3613, w3709};
	assign w1989 = w1508 ? w1988 : w1981;
	assign w1453 = w1451 & w1452;
	assign w1351 = {w1349, w1348};
	assign w101 = {w51, w100};
	assign w1456 = w1247;
	assign w1458 = w1240;
	assign w2307 = {w2306, w2305};
	assign w642 = w625 & w606;
	assign w1459 = w1297;
	assign w4373 = w4372 ? w3726 : s1780;
	assign w2603 = s2601;
	assign w1460 = w1238;
	assign w2486 = {w2485, w2484};
	assign w1461 = w1328;
	assign w2727 = w770;
	assign w1463 = i9;
	assign w4670 = w4669 & w3756;
	assign w1471 = w835 ? w1183 : w47;
	assign w4781 = w4780 ? w3726 : s1979;
	assign w4122 = w3770 & w4113;
	assign w1472 = w1183 ^ w1172;
	assign w316 = w308 != w44;
	assign w1324 = w1323;
	assign w1775 = w1499 ? w1774 : w1771;
	assign w4602 = w4601 ? w3726 : s1892;
	assign w1474 = w1473;
	assign w1477 = w829 ? w1476 : i25;
	assign w1478 = s1467[63:32];
	assign w1010 = s1009 & w1005;
	assign w103 = w102 ? w23 : w47;
	assign w1479 = {w832, w826};
	assign w2268 = i6[23:23];
	assign w1230 = i13;
	assign w1487 = w1244;
	assign w1489 = w788;
	assign w1705 = w1494 ? s1704 : s1703;
	assign w1494 = s1492[0:0];
	assign w3663 = {w1244, w47};
	assign w2322 = i6[15:15];
	assign w2463 = i6[15:15];
	assign w1495 = w1494 ? s1491 : s1490;
	assign w1972 = w1499 ? w1971 : w1968;
	assign w1473 = w826 ? w1472 : w1471;
	assign w1498 = w1494 ? s1497 : s1496;
	assign w2521 = w2502 ? w696 : i36;
	assign w80 = w27 & s55;
	assign w1580 = w1494 ? s1579 : s1578;
	assign w2348 = i6[15:15];
	assign w3631 = w3630 ? w367 : w3628;
	assign w3227 = s2760 == w3226;
	assign w780 = {w779, i1};
	assign w1503 = w1494 ? s1502 : s1501;
	assign w1506 = w1494 ? s1505 : s1504;
	assign w4863 = i13 ? w4862 : w47;
	assign w4773 = w4772 ? w3726 : s1976;
	assign w1508 = s1492[2:2];
	assign w3878 = w3877 & w3756;
	assign w204 = {2'b00, w203};
	assign w1388 = w1297[33:33];
	assign w1509 = w1508 ? w1507 : w1500;
	assign w4119 = w4118 & w3756;
	assign w3288 = i12 ? w3287 : w403;
	assign w2379 = i6[7:7];
	assign w1516 = w1499 ? w1515 : w1512;
	assign w1519 = w1494 ? s1518 : s1517;
	assign w2212 = {w2211, w2210};
	assign w4979 = i13 ? w4978 : w117;
	assign w2400 = {w2399, w2398};
	assign w4487 = w4486 ? w3726 : s1836;
	assign w229 = {w214, w228};
	assign w1525 = s1492[3:3];
	assign w1529 = w1494 ? s1528 : s1527;
	assign w1533 = w1499 ? w1532 : w1529;
	assign w3517 = w2706 ? w3516 : s813;
	assign w2833 = s305[31:31];
	assign w1883 = w1494 ? s1882 : s1881;
	assign w1536 = w1494 ? s1535 : s1534;
	assign w1957 = w1499 ? w1956 : w1953;
	assign w1540 = w1499 ? w1539 : w1536;
	assign w4913 = w3251 ? w4912 : w4909;
	assign w1334 = w1328[33:33];
	assign w1702 = w1508 ? w1701 : w1694;
	assign w1541 = w1508 ? w1540 : w1533;
	assign w1548 = w1499 ? w1547 : w1544;
	assign w1551 = w1494 ? s1550 : s1549;
	assign w1556 = w1508 ? w1555 : w1548;
	assign w4410 = w4409 ? w3726 : s1800;
	assign w1269 = w1268 ? w1267 : i24;
	assign w2738 = w913;
	assign w1559 = w1558 ? w1557 : w1526;
	assign w1562 = w1494 ? s1561 : s1560;
	assign w1565 = w1494 ? s1564 : s1563;
	assign w1569 = w1494 ? s1568 : s1567;
	assign w2105 = w2066;
	assign w1573 = w1499 ? w1572 : w1569;
	assign w2171 = w2020;
	assign w3374 = w3373 ? w3293 : s441;
	assign w1574 = w1508 ? w1573 : w1566;
	assign w1584 = w1494 ? s1583 : s1582;
	assign w1470 = s762;
	assign w2660 = 11'b11000110001;
	assign w1588 = w1499 ? w1587 : w1584;
	assign w1589 = w1508 ? w1588 : w1581;
	assign w1590 = w1525 ? w1589 : w1574;
	assign w558 = ~w557;
	assign w2328 = i6[15:15];
	assign w3142 = w398[2:2];
	assign w703 = s305[6:0];
	assign w915 = w736;
	assign w1593 = w1494 ? s1592 : s1591;
	assign w3409 = w3408 & w3313;
	assign w1310 = w1289[1:1];
	assign w2448 = {w2447, w2446};
	assign w200 = 10'b1100110011;
	assign w1596 = w1494 ? s1595 : s1594;
	assign w1090 = s18;
	assign w1597 = w1499 ? w1596 : w1593;
	assign w2032 = w2031 ? w2014 : w2029;
	assign w3491 = w3467 ? w3490 : w3487;
	assign w2643 = ~w2642;
	assign w1600 = w1494 ? s1599 : s1598;
	assign w4929 = s18 & w944;
	assign w1637 = w1494 ? s1636 : s1635;
	assign w1604 = w1499 ? w1603 : w1600;
	assign w1611 = w1494 ? s1610 : s1609;
	assign w1612 = w1499 ? w1611 : w1608;
	assign w4966 = w3243 ? w4965 : w4958;
	assign w1615 = w1494 ? s1614 : s1613;
	assign w2788 = {w2787, w2786};
	assign w1619 = w1499 ? w1618 : w1615;
	assign w1020 = s127 == w1019;
	assign w1624 = w1623 ? w1622 : w1559;
	assign w2300 = i6[23:16];
	assign w1627 = w1494 ? s1626 : s1625;
	assign w1798 = w1499 ? w1797 : w1794;
	assign w1645 = w1494 ? s1644 : s1643;
	assign w1642 = w1494 ? s1641 : s1640;
	assign w2584 = w59 ? w2583 : w2573;
	assign w1655 = w1525 ? w1654 : w1639;
	assign w2954 = {w2953, w2952};
	assign w2126 = w2013[29:20];
	assign w3791 = w3790 ? w3726 : s1502;
	assign w2165 = w2087;
	assign w1670 = w1508 ? w1669 : w1662;
	assign w2669 = 9'b000010000;
	assign w3705 = w3684 == w3704;
	assign w1673 = w1494 ? s1672 : s1671;
	assign w2244 = ~w741;
	assign w3310 = w3304 & w3309;
	assign w1680 = w1494 ? s1679 : s1678;
	assign w2147 = w2046;
	assign w1684 = w1499 ? w1683 : w1680;
	assign w1909 = w1499 ? w1908 : w1905;
	assign w1686 = w1525 ? w1685 : w1670;
	assign w3728 = {w47, s792};
	assign w2073 = w2013[31:20];
	assign w4192 = w4191 & w3756;
	assign w1464 = s127;
	assign w539 = ~w538;
	assign w1687 = w1558 ? w1686 : w1655;
	assign w4879 = s2626 + w4878;
	assign w1700 = w1494 ? s1699 : s1698;
	assign w1701 = w1499 ? w1700 : w1697;
	assign w1708 = w1494 ? s1707 : s1706;
	assign w4132 = w4131 ? w3726 : s1663;
	assign w1709 = w1499 ? w1708 : w1705;
	assign w3694 = {w3692, w3693};
	assign w1057 = {20'b00000000000000000000, w1056};
	assign w1712 = w1494 ? s1711 : s1710;
	assign w2277 = {w2276, w2275};
	assign w1431 = w1297[33:33];
	assign w1715 = w1494 ? s1714 : s1713;
	assign w1721 = w1494 ? s1720 : s1719;
	assign w1724 = w1494 ? s1723 : s1722;
	assign w1987 = w1494 ? s1986 : s1985;
	assign w1725 = w1499 ? w1724 : w1721;
	assign w1728 = w1494 ? s1727 : s1726;
	assign w2219 = i6[31:31];
	assign w1731 = w1494 ? s1730 : s1729;
	assign w4341 = w4340 ? w3726 : s1765;
	assign w1732 = w1499 ? w1731 : w1728;
	assign w2442 = {w2441, w2440};
	assign w1740 = w1499 ? w1739 : w1736;
	assign w3426 = w3302 & w3425;
	assign w2323 = {w2322, w2321};
	assign w1743 = w1494 ? s1742 : s1741;
	assign w2458 = {w2457, w2456};
	assign w1746 = w1494 ? s1745 : s1744;
	assign w3735 = w3734 == w47;
	assign w3539 = i13 ? w3538 : w47;
	assign w1747 = w1499 ? w1746 : w1743;
	assign w2396 = {w2395, w2394};
	assign w1748 = w1508 ? w1747 : w1740;
	assign w1756 = w1494 ? s1755 : s1754;
	assign w3763 = w3762 & w3753;
	assign w1760 = w1499 ? w1759 : w1756;
	assign w1763 = w1494 ? s1762 : s1761;
	assign w3682 = s1294[34:34];
	assign w801 = ~w800;
	assign w1771 = w1494 ? s1770 : s1769;
	assign w3639 = w3638 == w34;
	assign w1778 = w1494 ? s1777 : s1776;
	assign w3211 = {w3195, w3191};
	assign w1781 = w1494 ? s1780 : s1779;
	assign w4947 = s2999[31:1];
	assign w1783 = w1508 ? w1782 : w1775;
	assign w2365 = i6[7:7];
	assign w1784 = w1525 ? w1783 : w1768;
	assign w1790 = w1494 ? s1789 : s1788;
	assign w2378 = {w2377, w2376};
	assign w1791 = w1499 ? w1790 : w1787;
	assign w1802 = w1494 ? s1801 : s1800;
	assign w962 = {w186, w183};
	assign w1805 = w1494 ? s1804 : s1803;
	assign w1355 = w1328[33:33];
	assign w1806 = w1499 ? w1805 : w1802;
	assign w2213 = i6[31:31];
	assign w3166 = w3142 ? w3165 : w3162;
	assign w1323 = -w1322;
	assign w1812 = w1494 ? s1811 : s1810;
	assign w362 = w311 == w361;
	assign w1908 = w1494 ? s1907 : s1906;
	assign w2242 = w741 ? w2241 : i28;
	assign w3945 = w3944 & w3756;
	assign w2194 = {w2193, w2192};
	assign w687 = 12'b111111111111;
	assign w2382 = {w2381, w2380};
	assign w1814 = w1508 ? w1813 : w1806;
	assign w1739 = w1494 ? s1738 : s1737;
	assign w1819 = w1494 ? s1818 : s1817;
	assign w971 = {1'b0, w23};
	assign w315 = w314 ? w310 : w301;
	assign w1822 = w1494 ? s1821 : s1820;
	assign w161 = {4'b0000, w160};
	assign w1823 = w1499 ? w1822 : w1819;
	assign w2734 = w982;
	assign w1829 = w1494 ? s1828 : s1827;
	assign w4811 = w3820 & w4766;
	assign w3855 = w3854 ? w3726 : s1528;
	assign w800 = w796 == w799;
	assign w1830 = w1499 ? w1829 : w1826;
	assign w1831 = w1508 ? w1830 : w1823;
	assign w2297 = {w2296, w2295};
	assign w4542 = w3810 & w4505;
	assign w1834 = w1494 ? s1833 : s1832;
	assign w1837 = w1494 ? s1836 : s1835;
	assign w1838 = w1499 ? w1837 : w1834;
	assign w838 = {w835, w837};
	assign w1844 = w1494 ? s1843 : s1842;
	assign w376 = w375 ? w367 : w366;
	assign w1845 = w1499 ? w1844 : w1841;
	assign w1846 = w1508 ? w1845 : w1838;
	assign w740 = w736[9:9];
	assign w2822 = w337 ? w2821 : w2820;
	assign w3261 = s235[0:0];
	assign w1847 = w1525 ? w1846 : w1831;
	assign w1850 = w1494 ? s1849 : s1848;
	assign w482 = {s475, w481};
	assign w1853 = w1494 ? s1852 : s1851;
	assign w3838 = w3837 & w3756;
	assign w2570 = {w23, w2569};
	assign w1861 = w1499 ? w1860 : w1857;
	assign w1865 = w1494 ? s1864 : s1863;
	assign w1352 = w1328[33:33];
	assign w1925 = w1499 ? w1924 : w1921;
	assign w4070 = w4069 & w3756;
	assign w1869 = w1499 ? w1868 : w1865;
	assign w507 = w484[191:160];
	assign w2340 = i6[15:15];
	assign w1878 = w1525 ? w1877 : w1862;
	assign w1880 = w1623 ? w1879 : w1816;
	assign w3259 = i12 ? w3258 : s180;
	assign w296 = w240 | w295;
	assign w1895 = w1508 ? w1894 : w1887;
	assign w3687 = ~w3686;
	assign w1898 = w1494 ? s1897 : s1896;
	assign w3875 = w3874 ? w3726 : s1537;
	assign w2761 = w737;
	assign w1901 = w1494 ? s1900 : s1899;
	assign w1902 = w1499 ? w1901 : w1898;
	assign w1914 = w1494 ? s1913 : s1912;
	assign w4215 = w3810 & w4178;
	assign w3700 = s1294[17:1];
	assign w2107 = w788;
	assign w1921 = w1494 ? s1920 : s1919;
	assign w3461 = w3459 ? s418 : s417;
	assign w136 = 6'b110111;
	assign w2106 = w2076;
	assign w1929 = w1494 ? s1928 : s1927;
	assign w2180 = w61;
	assign w1933 = w1499 ? w1932 : w1929;
	assign w4023 = w4022 & w3756;
	assign w1939 = w1494 ? s1938 : s1937;
	assign w1940 = w1499 ? w1939 : w1936;
	assign w4977 = w3243 ? w4976 : w4974;
	assign w540 = w539 | w493;
	assign w1941 = w1508 ? w1940 : w1933;
	assign w4134 = w3788 & w4113;
	assign w1958 = w1508 ? w1957 : w1950;
	assign w1964 = w1494 ? s1963 : s1962;
	assign w2656 = {2'b00, w2655};
	assign w2202 = {w2201, w2200};
	assign w1974 = w1525 ? w1973 : w1958;
	assign w4298 = w4297 ? w3726 : s1742;
	assign w2403 = i6[7:7];
	assign w4345 = w4344 ? w3726 : s1769;
	assign w1981 = w1499 ? w1980 : w1977;
	assign w1971 = w1494 ? s1970 : s1969;
	assign w2225 = i6[31:31];
	assign w4343 = w3805 & w4310;
	assign w3015 = w946;
	assign w2419 = i6[31:31];
	assign w1330 = {w1328, w403};
	assign w1984 = w1494 ? s1983 : s1982;
	assign w1587 = w1494 ? s1586 : s1585;
	assign w1618 = w1494 ? s1617 : s1616;
	assign w1995 = w1494 ? s1994 : s1993;
	assign w1996 = w1499 ? w1995 : w1992;
	assign w2002 = w1494 ? s2001 : s2000;
	assign w2158 = w2014;
	assign w2003 = w1499 ? w2002 : w1999;
	assign w3772 = w3771 & w3756;
	assign w2804 = s305[31:31];
	assign w607 = w551 & w606;
	assign w2005 = w1525 ? w2004 : w1989;
	assign w2007 = w1623 ? w2006 : w1943;
	assign w4166 = w3831 & w4113;
	assign w3401 = w3400 ? w3293 : s455;
	assign w479 = {s472, w478};
	assign w2009 = w47 ? w2008 : w1753;
	assign w724 = {w47, w723};
	assign w2647 = 9'b000000000;
	assign w1364 = w1328[33:33];
	assign w2010 = w808 ? w2009 : w303;
	assign w2011 = 31'b0000000000000000000000000000000;
	assign w2012 = {w2011, i1};
	assign w4024 = w4023 ? w3726 : s1609;
	assign w1064 = w1063 ? w1060 : w1059;
	assign w2014 = w2013[24:20];
	assign w2015 = w2014;
	assign w2018 = w2013[19:15];
	assign w2021 = w2020;
	assign w2024 = {w23, w2023};
	assign w2027 = w2026 ? w2018 : w2024;
	assign w2677 = w2649 == w2676;
	assign w3293 = i12 ? w3292 : i38;
	assign w2029 = {w23, w2028};
	assign w2631 = s2615;
	assign w2030 = |w2014;
	assign w2876 = {w2875, w2874};
	assign w918 = {w156, w186};
	assign w32 = 2'b10;
	assign w2427 = i6[31:31];
	assign w3832 = w3831 & w3753;
	assign w3468 = w3467 ? w3466 : w3463;
	assign w3371 = w3334 & w3353;
	assign w2031 = ~w2030;
	assign w2036 = {w2027, w2034};
	assign w4730 = w3798 & w4701;
	assign w2038 = {w2032, w2036};
	assign w1295 = s1294[34:1];
	assign w2039 = w2013[29:25];
	assign w34 = 2'b11;
	assign w2043 = w2013[6:0];
	assign w195 = {3'b000, w194};
	assign w2047 = {1'b0, w32};
	assign w3905 = w3836 & w3848;
	assign w3165 = w3137 ? w3164 : w3163;
	assign w2897 = s305[31:31];
	assign w1753 = w1752 ? w1751 : w1624;
	assign w2369 = i6[7:7];
	assign w2052 = {w23, w2051};
	assign w4532 = w4531 ? w3726 : s1858;
	assign w2053 = |w2020;
	assign w2054 = ~w2053;
	assign w3953 = w3952 & w3756;
	assign w2635 = w2634;
	assign w2057 = {w2055, w2056};
	assign w134 = s127 == w133;
	assign w2060 = {w2027, w2059};
	assign w179 = w178 ? s152 : w47;
	assign w2061 = w2013[29:20];
	assign w1653 = w1499 ? w1652 : w1649;
	assign w2062 = {w2061, w2060};
	assign w2063 = {w2033, w2062};
	assign w2065 = w2043 == w2064;
	assign w232 = {w219, w230};
	assign w2070 = w2013[14:12];
	assign w2071 = {w2070, w2069};
	assign w2079 = {w2055, w2078};
	assign w1222 = w1221;
	assign w2074 = {w2073, w2072};
	assign w2075 = {2'b00, w184};
	assign w2671 = {2'b00, w2670};
	assign w2076 = w2043 == w2075;
	assign w2082 = {w2027, w2081};
	assign w2460 = {w2459, w2458};
	assign w2083 = {w2032, w2082};
	assign w4743 = w4742 & w3756;
	assign w2084 = w2013[31:25];
	assign w1076 = s813;
	assign w2663 = w2662 ? w2659 : w2658;
	assign w4777 = w4776 ? w3726 : s1978;
	assign w2086 = {1'b0, w181};
	assign w4079 = w4078 ? w3726 : s1636;
	assign w1500 = w1499 ? w1498 : w1495;
	assign w2088 = w2087 ? w2085 : w2077;
	assign w1767 = w1499 ? w1766 : w1763;
	assign w2562 = w278 ? w2561 : w2560;
	assign w3941 = w3940 & w3756;
	assign w1926 = w1508 ? w1925 : w1918;
	assign w2089 = w2088;
	assign w2092 = w2013[31:25];
	assign w2094 = w2020;
	assign w2100 = i2;
	assign w1243 = {1'b0, w1242};
	assign w1652 = w1494 ? s1651 : s1650;
	assign w2101 = w23;
	assign w2102 = i9;
	assign w2103 = w2049;
	assign w1271 = s1270 == w544;
	assign w2108 = i9;
	assign w4859 = w4858 ? w47 : w4855;
	assign w3707 = w1312 ? w3706 : s1294;
	assign w695 = w316 ? w692 : w687;
	assign w60 = w59 ? w57 : w52;
	assign w2708 = w2692[2:2];
	assign w2109 = w808;
	assign w2264 = i6[23:23];
	assign w2110 = i2;
	assign w4535 = w4534 & w3756;
	assign w600 = w597 | w599;
	assign w2383 = i6[7:7];
	assign w2116 = w781;
	assign w2536 = w45;
	assign w2404 = {w2403, w2402};
	assign w2117 = w2013;
	assign w2118 = w775;
	assign w2646 = s896;
	assign w2120 = w2074;
	assign w3783 = w3736 & w3782;
	assign w2546 = i5 ? w696 : w86;
	assign w2122 = {w2055, w2121};
	assign w2125 = {w2027, w2124};
	assign w2128 = w2127;
	assign w1862 = w1508 ? w1861 : w1854;
	assign w2130 = w2013[14:0];
	assign w2935 = s305[31:31];
	assign w2131 = {w2027, w2130};
	assign w43 = w29 ? w42 : i15;
	assign w2132 = {w2032, w2131};
	assign w2757 = w811;
	assign w2135 = w2134;
	assign w4887 = w2716 ? w23 : w47;
	assign w1327 = w1238 + w1323;
	assign w2136 = w2076;
	assign w1115 = i12;
	assign w2214 = {w2213, w2212};
	assign w2139 = w2049;
	assign w2940 = {w2939, w2938};
	assign w2141 = w2140;
	assign w2695 = w2694;
	assign w201 = {2'b00, w200};
	assign w2640 = i9;
	assign w2143 = w2142;
	assign w2146 = w2032;
	assign w1062 = {20'b00000000000000000000, w1061};
	assign w2148 = w2092;
	assign w2151 = w2092;
	assign w1309 = w1308;
	assign w2389 = i6[7:7];
	assign w2152 = w2043;
	assign w845 = s127 == w844;
	assign w2155 = w2020;
	assign w2156 = w2018;
	assign w2983 = i13;
	assign w2355 = {w2353, w2354};
	assign w2157 = w2014;
	assign w3590 = w3589 == w34;
	assign w2159 = w23;
	assign w4470 = w4469 & w3756;
	assign w2162 = w2088;
	assign w2164 = w2066;
	assign w585 = w584 & w558;
	assign w2166 = w2049;
	assign w2096 = w2095;
	assign w2167 = w2046;
	assign w2168 = w2092;
	assign w2169 = w2013;
	assign w2170 = w2095;
	assign w1114 = w770;
	assign w2172 = w2092;
	assign w2332 = i6[15:15];
	assign w2391 = i6[7:7];
	assign w156 = s127 == w155;
	assign w2692 = w2691 ? w2689 : w2688;
	assign w3610 = w3589 == w3609;
	assign w2174 = w2020;
	assign w2945 = s305[31:31];
	assign w2175 = w2018;
	assign w2176 = w2014;
	assign w2557 = {w47, w2556};
	assign w3836 = w3769 & w3825;
	assign w2209 = i6[31:31];
	assign w2844 = {w2843, w2842};
	assign w3991 = w3990 & w3756;
	assign w1466 = w770;
	assign w2177 = w2014;
	assign w2178 = w38;
	assign w2179 = i3;
	assign w2182 = i4;
	assign w2184 = w97;
	assign w2471 = i6[15:15];
	assign w2186 = w105;
	assign w1016 = w956 ? w1015 : w1014;
	assign w2616 = i13;
	assign w2198 = {w2197, w2196};
	assign w1029 = w1028;
	assign w2231 = i6[31:31];
	assign w1425 = w1297[33:33];
	assign w2199 = i6[31:31];
	assign w2200 = {w2199, w2198};
	assign w2342 = i6[15:15];
	assign w2203 = i6[31:31];
	assign w4654 = w4653 & w3756;
	assign w2204 = {w2203, w2202};
	assign w1113 = i9;
	assign w2206 = {w2205, w2204};
	assign w811 = w810 ? w47 : w23;
	assign w2207 = i6[31:31];
	assign w2566 = w100 ? w2565 : w2563;
	assign w2210 = {w2209, w2208};
	assign w2215 = i6[31:31];
	assign w3776 = w3775 & w3741;
	assign w717 = s305[6:0];
	assign w2510 = {w2509, w2508};
	assign w2887 = s305[31:31];
	assign w2220 = {w2219, w2218};
	assign w2299 = w2244 ? w2243 : w2298;
	assign w4577 = w4576 & w3756;
	assign w1961 = w1494 ? s1960 : s1959;
	assign w2490 = ~w2452;
	assign w398 = w299 ? w397 : w376;
	assign w2223 = i6[31:31];
	assign w2226 = {w2225, w2224};
	assign w3665 = w1259 ? w3664 : w3661;
	assign w2193 = i6[31:31];
	assign w2227 = i6[31:31];
	assign w225 = {w202, w224};
	assign w2229 = i6[31:31];
	assign w143 = 7'b1110011;
	assign w2706 = w2692[8:8];
	assign w689 = s305[6:0];
	assign w2230 = {w2229, w2228};
	assign w2233 = {w2231, w2230};
	assign w2234 = i6[31:31];
	assign w2236 = {w2234, w2233};
	assign w2239 = {w2237, w2236};
	assign w2240 = i6[31:31];
	assign w3344 = w3324 & w3335;
	assign w3196 = w3195 ? w3193 : w3192;
	assign w2352 = w741 ? w2351 : i30;
	assign w3395 = w3318 & w3390;
	assign w2245 = w2244 ? w2243 : w2242;
	assign w2563 = w76 ? w2562 : w2555;
	assign w2993 = i13;
	assign w2246 = i6[31:24];
	assign w2249 = w2248 ? w2247 : i27;
	assign w2251 = i6[23:23];
	assign w2255 = {w2254, w2253};
	assign w2823 = w340 ? w2812 : w2822;
	assign w2257 = {w2256, w2255};
	assign w1143 = w1130 ? w23 : w47;
	assign w2258 = i6[23:23];
	assign w2262 = i6[23:23];
	assign w2265 = {w2264, w2263};
	assign w2811 = s305[31:31];
	assign w2864 = {w2863, w2862};
	assign w2019 = w2018;
	assign w2267 = {w2266, w2265};
	assign w2269 = {w2268, w2267};
	assign w4359 = w3826 & w4310;
	assign w2008 = w1752 ? w2007 : w1880;
	assign w2270 = i6[23:23];
	assign w2318 = i6[15:15];
	assign w2273 = {w2272, w2271};
	assign w2274 = i6[23:23];
	assign w2278 = i6[23:23];
	assign w4454 = w4453 & w3756;
	assign w1558 = s1492[4:4];
	assign w2279 = {w2278, w2277};
	assign w4250 = w4249 ? w3726 : s1720;
	assign w2506 = {w2505, w2504};
	assign w2736 = i9;
	assign w2281 = {w2280, w2279};
	assign w1936 = w1494 ? s1935 : s1934;
	assign w2282 = i6[23:23];
	assign w2741 = w890;
	assign w2351 = {w2350, w2349};
	assign w2284 = i6[23:23];
	assign w1058 = s19 == w1057;
	assign w2285 = {w2284, w2283};
	assign w2371 = i6[7:7];
	assign w2286 = i6[23:23];
	assign w4225 = w4224 ? w3726 : s1707;
	assign w2287 = {w2286, w2285};
	assign w1876 = w1499 ? w1875 : w1872;
	assign w2511 = w2413 ? w2510 : w117;
	assign w2288 = i6[23:23];
	assign w4339 = w3798 & w4310;
	assign w2289 = {w2288, w2287};
	assign w1188 = w1187[31:16];
	assign w2291 = {w2290, w2289};
	assign w4719 = w4718 & w3756;
	assign w2292 = i6[23:23];
	assign w2728 = w770;
	assign w1768 = w1508 ? w1767 : w1760;
	assign w2293 = {w2292, w2291};
	assign w2295 = {w2294, w2293};
	assign w3049 = {w199, w193};
	assign w2296 = i6[23:23];
	assign w2298 = w741 ? w2297 : i29;
	assign w2301 = {w2299, w2300};
	assign w4984 = s18 ^ w944;
	assign w2303 = w2302 ? w2301 : w2249;
	assign w2305 = i6[15:15];
	assign w4441 = w3742 & w4440;
	assign w3976 = w3841 & w3915;
	assign w2408 = w2244 ? w2243 : w2407;
	assign w2306 = i6[15:15];
	assign w3674 = s1270 + w3673;
	assign w2308 = i6[15:15];
	assign w3706 = w3705 ? w3703 : w3698;
	assign w3218 = i13 ? w2517 : w117;
	assign w2310 = i6[15:15];
	assign w2376 = {w2375, w2374};
	assign w2312 = i6[15:15];
	assign w188 = 9'b110110011;
	assign w1361 = w1328[33:33];
	assign w2313 = {w2312, w2311};
	assign w3024 = w3023 ? s3000 : i37;
	assign w2319 = {w2318, w2317};
	assign w529 = s444 == s475;
	assign w2320 = i6[15:15];
	assign w2325 = {w2324, w2323};
	assign w2681 = {3'b000, w2680};
	assign w2326 = i6[15:15];
	assign w2327 = {w2326, w2325};
	assign w778 = w776 & w777;
	assign w1946 = w1494 ? s1945 : s1944;
	assign w2447 = i6[31:31];
	assign w2329 = {w2328, w2327};
	assign w2330 = i6[15:15];
	assign w4027 = w4026 & w3756;
	assign w2331 = {w2330, w2329};
	assign w481 = {s474, w480};
	assign w2333 = {w2332, w2331};
	assign w2893 = s305[31:31];
	assign w2334 = i6[15:15];
	assign w2335 = {w2334, w2333};
	assign w3994 = w3776 & w3981;
	assign w738 = w737;
	assign w933 = {w183, w932};
	assign w396 = w319 ? w377 : w301;
	assign w2336 = i6[15:15];
	assign w2712 = w2692[5:5];
	assign w483 = w47 ? w482 : w467;
	assign w2338 = i6[15:15];
	assign w65 = {w27, w25};
	assign w2341 = {w2340, w2339};
	assign w3873 = w3793 & w3848;
	assign w2436 = {w2435, w2434};
	assign w2343 = {w2342, w2341};
	assign w2345 = {w2344, w2343};
	assign w2349 = {w2348, w2347};
	assign w2350 = i6[15:15];
	assign w2353 = w2244 ? w2243 : w2352;
	assign w1430 = {w1429, w1428};
	assign w2357 = w974 == w2356;
	assign w2358 = w2357 ? w2355 : w2303;
	assign w3612 = w1198 ? w3611 : s1160;
	assign w1577 = w1494 ? s1576 : s1575;
	assign w2362 = {w2361, w2360};
	assign w2363 = i6[7:7];
	assign w4972 = s3001[30:0];
	assign w2364 = {w2363, w2362};
	assign w4031 = w4030 & w3756;
	assign w2366 = {w2365, w2364};
	assign w2137 = w2066;
	assign w2373 = i6[7:7];
	assign w2374 = {w2373, w2372};
	assign w3754 = w3742 & w3753;
	assign w2380 = {w2379, w2378};
	assign w2894 = {w2893, w2892};
	assign w2381 = i6[7:7];
	assign w3301 = w3300 == w47;
	assign w2755 = w2754;
	assign w2384 = {w2383, w2382};
	assign w2387 = i6[7:7];
	assign w2006 = w1558 ? w2005 : w1974;
	assign w2388 = {w2387, w2386};
	assign w2854 = {w2853, w2852};
	assign w476 = {s469, s468};
	assign w2390 = {w2389, w2388};
	assign w519 = s439 == s470;
	assign w2774 = {w2773, w2772};
	assign w2392 = {w2391, w2390};
	assign w2393 = i6[7:7];
	assign w434 = {s421, w432};
	assign w2394 = {w2393, w2392};
	assign w2470 = {w2469, w2468};
	assign w2398 = {w2397, w2396};
	assign w2720 = w2693;
	assign w4576 = w3762 & w4571;
	assign w276 = w275 ? w23 : w273;
	assign w2405 = i6[7:7];
	assign w1256 = {17'b00000000000000000, w23};
	assign w851 = s127 == w850;
	assign w1877 = w1508 ? w1876 : w1869;
	assign w2195 = i6[31:31];
	assign w2406 = {w2405, w2404};
	assign w2407 = w741 ? w2406 : i31;
	assign w2409 = i6[7:0];
	assign w1067 = 32'b00000000000000000000000000000001;
	assign w2411 = w976 ? w2410 : w2358;
	assign w2412 = |w737;
	assign w1669 = w1499 ? w1668 : w1665;
	assign w2160 = i2;
	assign w2417 = w2244 ? w403 : i33;
	assign w859 = s127 == w858;
	assign w2418 = i6[31:31];
	assign w3778 = w3777 & w3756;
	assign w3250 = {2'b00, w32};
	assign w1749 = w1525 ? w1748 : w1733;
	assign w2421 = i6[31:31];
	assign w2827 = s305[31:31];
	assign w2422 = {w2421, w2420};
	assign w2423 = i6[31:31];
	assign w2426 = {w2425, w2424};
	assign w3867 = w3866 ? w3726 : s1534;
	assign w2522 = {3'b000, w23};
	assign w4205 = w4204 ? w3726 : s1698;
	assign w731 = w362 ? w730 : w729;
	assign w2428 = {w2427, w2426};
	assign w3209 = w3187 ? w47 : w3208;
	assign w1977 = w1494 ? s1976 : s1975;
	assign w2739 = w294;
	assign w843 = 10'b1111100011;
	assign w2430 = {w2429, w2428};
	assign w2080 = w2013[14:12];
	assign w2432 = {w2431, w2430};
	assign w3129 = w679;
	assign w2433 = i6[31:31];
	assign w4566 = w3841 & w4505;
	assign w3678 = w3677 ? w367 : w3675;
	assign w741 = ~w740;
	assign w2747 = w2746;
	assign w4953 = s2995 ? w4952 : s18;
	assign w2437 = i6[31:31];
	assign w2438 = {w2437, w2436};
	assign w1337 = w1328[33:33];
	assign w2440 = {w2439, w2438};
	assign w3031 = {w848, w845};
	assign w2443 = i6[31:31];
	assign w145 = s127 == w144;
	assign w2444 = {w2443, w2442};
	assign w3906 = w3905 & w3756;
	assign w2445 = i6[31:31];
	assign w3473 = w3459 ? s444 : s443;
	assign w2539 = i9;
	assign w168 = {2'b00, w167};
	assign w2449 = w741 ? w2448 : w2417;
	assign w2452 = w20[1:1];
	assign w1248 = {1'b0, w1247};
	assign w2455 = w2244 ? w403 : i34;
	assign w2457 = i6[15:15];
	assign w2866 = {w2865, w2864};
	assign w2461 = i6[15:15];
	assign w4349 = w4348 ? w3726 : s1770;
	assign w2718 = w2692[4:4];
	assign w2549 = {w47, w2548};
	assign w2464 = {w2463, w2462};
	assign w568 = w567 & w562;
	assign w2466 = {w2465, w2464};
	assign w4918 = 4'b0001;
	assign w2468 = {w2467, w2466};
	assign w349 = w348 ? w345 : w341;
	assign w25 = s22 == w24;
	assign w2852 = {w2851, w2850};
	assign w875 = {w208, w873};
	assign w2472 = {w2471, w2470};
	assign w2474 = {w2473, w2472};
	assign w2475 = i6[15:15];
	assign w2476 = {w2475, w2474};
	assign w3599 = {w3597, w3598};
	assign w2477 = i6[15:15];
	assign w4572 = w3742 & w4571;
	assign w2480 = {w2479, w2478};
	assign w3932 = w3783 & w3915;
	assign w2629 = s2596;
	assign w2483 = i6[15:15];
	assign w2484 = {w2483, w2482};
	assign w2485 = i6[15:15];
	assign w2487 = w741 ? w2486 : w2455;
	assign w3444 = w3443 & w3313;
	assign w2489 = {w2487, w2488};
	assign w2493 = w979 ? i6 : w2492;
	assign w2496 = w2495;
	assign w2793 = s305[31:31];
	assign w2498 = s22;
	assign w2500 = {w33, w25};
	assign w28 = {w27, w25};
	assign w716 = {w715, w714};
	assign w2501 = {w35, w2500};
	assign w2502 = |w2501;
	assign w2119 = w811;
	assign w2504 = s762[7:0];
	assign w2221 = i6[31:31];
	assign w2505 = s762[7:0];
	assign w2508 = {w2507, w2506};
	assign w1063 = s19 == w1062;
	assign w2512 = s762[15:0];
	assign w2513 = s762[15:0];
	assign w2795 = s305[31:31];
	assign w2517 = w27 ? w2516 : w2503;
	assign w2764 = w2763;
	assign w659 = ~w658;
	assign w2518 = w2517;
	assign w4813 = w4812 ? w3726 : s1994;
	assign w2809 = s305[31:31];
	assign w2523 = {2'b00, w974};
	assign w2271 = {w2270, w2269};
	assign w2526 = 4'b0011;
	assign w3703 = {w3702, w3701};
	assign w339 = {2'b00, w184};
	assign w2528 = w2452 ? w2527 : w2526;
	assign w622 = w584 & w612;
	assign w2435 = i6[31:31];
	assign w2529 = w972 ? w2528 : w2525;
	assign w2530 = 4'b1111;
	assign w1046 = 12'b110000000001;
	assign w2532 = w27 ? w2531 : w2521;
	assign w4034 = w3831 & w3981;
	assign w3995 = w3994 & w3756;
	assign w748 = w319 ? w367 : w747;
	assign w2824 = s305[11:7];
	assign w4246 = w4245 ? w3726 : s1719;
	assign w850 = {2'b00, w849};
	assign w2534 = w115;
	assign w2535 = w982;
	assign w2537 = w69;
	assign w2540 = w294;
	assign w2542 = w249;
	assign w827 = 11'b10000110011;
	assign w2545 = s305;
	assign w2791 = s305[31:31];
	assign w730 = w359 ? w692 : w687;
	assign w1816 = w1558 ? w1815 : w1784;
	assign w2547 = w87 ? w2546 : w696;
	assign w374 = {w372, w373};
	assign w2548 = w258 ? w42 : w71;
	assign w2553 = {w47, w2552};
	assign w2798 = s305[31:31];
	assign w4907 = w3187 ? w2561 : w4906;
	assign w2556 = w270 ? w42 : w74;
	assign w944 = w943 ? s762 : w927;
	assign w2559 = 4'b0111;
	assign w2564 = i7 ? w688 : w34;
	assign w2561 = 4'b0110;
	assign w4103 = w4102 ? w3726 : s1648;
	assign w2569 = w2568 ? w23 : w47;
	assign w1485 = w1251;
	assign w2571 = w244 ? w688 : w2570;
	assign w2574 = w272 ? w86 : s49;
	assign w319 = ~w318;
	assign w2625 = s2624 & w1067;
	assign w799 = {1'b0, s797};
	assign w2575 = w275 ? w2559 : w2574;
	assign w1204 = w1130 ? w34 : w688;
	assign w1774 = w1494 ? s1773 : s1772;
	assign w2580 = 3'b001;
	assign w2581 = {w2580, w2569};
	assign w2585 = w2584;
	assign w4710 = w3770 & w4701;
	assign w1766 = w1494 ? s1765 : s1764;
	assign w1736 = w1494 ? s1735 : s1734;
	assign w2599 = s2597;
	assign w2608 = i9;
	assign w2613 = s2612 ? s2611 : w47;
	assign w2399 = i6[7:7];
	assign w2620 = s2618;
	assign w564 = 6'b100000;
	assign w289 = w288 ? w23 : w287;
	assign w2622 = i13;
	assign w2957 = w2956 ? w2954 : w2951;
	assign w2628 = s2600;
	assign w1155 = w1130;
	assign w2636 = s984;
	assign w4015 = w4014 & w3756;
	assign w2488 = i6[15:0];
	assign w2642 = s18 | s19;
	assign w2594 = w741;
	assign w2644 = w2643 & s2632;
	assign w2648 = 9'b100000000;
	assign w2649 = {s127, w47};
	assign w2655 = 11'b11100110001;
	assign w4380 = w3762 & w4375;
	assign w504 = w488[159:128];
	assign w2661 = {2'b00, w2660};
	assign w4364 = w4363 & w3756;
	assign w2664 = 9'b000100000;
	assign w451 = {s444, w450};
	assign w2665 = 11'b10100110001;
	assign w2478 = {w2477, w2476};
	assign w2666 = {2'b00, w2665};
	assign w2667 = w2649 == w2666;
	assign w2668 = w2667 ? w2664 : w2663;
	assign w4035 = w4034 & w3756;
	assign w2670 = 11'b10000110001;
	assign w3287 = s409 + w3286;
	assign w978 = s55 ? w977 : w23;
	assign w2674 = 9'b000001000;
	assign w3666 = i13 ? w3665 : w3633;
	assign w2577 = 4'b0101;
	assign w2676 = {3'b000, w2675};
	assign w2678 = w2677 ? w2674 : w2673;
	assign w2784 = {w2783, w2782};
	assign w4285 = w4284 & w3756;
	assign w2679 = 9'b000000100;
	assign w1634 = w1494 ? s1633 : s1632;
	assign w2818 = w316 ? w2817 : w2767;
	assign w684 = ~w23;
	assign w2680 = 10'b1000110001;
	assign w4596 = w3793 & w4571;
	assign w4126 = w3776 & w4113;
	assign w3756 = w775 ? w47 : w3755;
	assign w2682 = w2649 == w2681;
	assign w1414 = {w1412, w1411};
	assign w2684 = 9'b000000010;
	assign w2685 = 9'b100110001;
	assign w2686 = {4'b0000, w2685};
	assign w2689 = 9'b000000001;
	assign w2697 = i10;
	assign w2699 = w2692;
	assign w502 = w498 & w501;
	assign w2707 = w2706;
	assign w2316 = i6[15:15];
	assign w2709 = w2708;
	assign w2710 = w2692[1:1];
	assign w1175 = w1174[31:16];
	assign w2713 = w2712;
	assign w4855 = w4854 ? w23 : w47;
	assign w3692 = w3691 + w1308;
	assign w523 = s441 == s472;
	assign w2716 = w2692[0:0];
	assign w2645 = w2644;
	assign w2717 = w2716;
	assign w2719 = w2718;
	assign w2721 = w2692[3:3];
	assign w2725 = s815;
	assign w2337 = {w2336, w2335};
	assign w2754 = w2753 ? w23 : w47;
	assign w2731 = s762;
	assign w3284 = i12 ? w3283 : w403;
	assign w2735 = w293;
	assign w2792 = {w2791, w2790};
	assign w2742 = &w736;
	assign w2967 = s18;
	assign w2744 = {4'b0000, w2743};
	assign w3934 = w3933 ? w3726 : s1567;
	assign w2746 = w2742 | w2745;
	assign w2503 = w2502 ? w117 : i35;
	assign w2748 = w736[6:0];
	assign w3548 = w2712 ? w117 : s984;
	assign w2750 = w2748 == w2749;
	assign w3800 = w3799 & w3756;
	assign w2753 = w2750 | w2752;
	assign w3255 = s2760 == w3254;
	assign w256 = i5 ? w47 : w23;
	assign w2756 = i12;
	assign w2759 = w741;
	assign w1315 = s180;
	assign w2762 = w736[5:5];
	assign w2763 = ~w2762;
	assign w3484 = w3467 ? w3483 : w3480;
	assign w2765 = i9;
	assign w4772 = w4771 & w3756;
	assign w4042 = w3841 & w3981;
	assign w2767 = 32'b11111111111111111111111111111111;
	assign w2832 = {w2831, w2830};
	assign w2769 = s305[31:31];
	assign w3907 = w3906 ? w3726 : s1552;
	assign w2770 = {w2769, w2768};
	assign w2771 = s305[31:31];
	assign w2772 = {w2771, w2770};
	assign w2020 = w2013[11:7];
	assign w2778 = {w2777, w2776};
	assign w2779 = s305[31:31];
	assign w3053 = |w3052;
	assign w1572 = w1494 ? s1571 : s1570;
	assign w2781 = s305[31:31];
	assign w2783 = s305[31:31];
	assign w2785 = s305[31:31];
	assign w2787 = s305[31:31];
	assign w4974 = w3240 ? w4973 : s3001;
	assign w4061 = w3776 & w4048;
	assign w2790 = {w2789, w2788};
	assign w2794 = {w2793, w2792};
	assign w4376 = w3742 & w4375;
	assign w4039 = w4038 & w3756;
	assign w148 = {w142, w147};
	assign w2797 = {w2795, w2794};
	assign w2800 = {w2798, w2797};
	assign w4755 = w4754 & w3756;
	assign w2803 = {w2801, w2800};
	assign w2806 = {w2804, w2803};
	assign w2807 = s305[31:31];
	assign w2808 = {w2807, w2806};
	assign w2810 = {w2809, w2808};
	assign w2812 = {w2811, w2810};
	assign w3192 = w3191 ? w3189 : w3182;
	assign w2814 = w314 ? w2813 : w2767;
	assign w3527 = w2694 ? w47 : s896;
	assign w2254 = i6[23:23];
	assign w2816 = s305[31:20];
	assign w3292 = w299 ? w770 : i39;
	assign w1272 = w1271 ? w23 : w47;
	assign w2819 = w319 ? w2817 : w2818;
	assign w331 = s305[14:14];
	assign w1630 = w1494 ? s1629 : s1628;
	assign w2820 = w321 ? w2819 : w2814;
	assign w2821 = w334 ? w117 : w2767;
	assign w2826 = {w2825, w2824};
	assign w1694 = w1499 ? w1693 : w1690;
	assign w2828 = {w2827, w2826};
	assign w2829 = s305[31:31];
	assign w804 = w776 & i2;
	assign w787 = w786 & w249;
	assign w2830 = {w2829, w2828};
	assign w2831 = s305[31:31];
	assign w4099 = w4098 ? w3726 : s1647;
	assign w2908 = {w2907, w2906};
	assign w2836 = {w2835, w2834};
	assign w2838 = {w2837, w2836};
	assign w2840 = {w2839, w2838};
	assign w4371 = w3841 & w4310;
	assign w2860 = {w2859, w2858};
	assign w2841 = s305[31:31];
	assign w2843 = s305[31:31];
	assign w2845 = s305[31:31];
	assign w2846 = {w2845, w2844};
	assign w3016 = w954;
	assign w2847 = s305[31:31];
	assign w2514 = {w2513, w2512};
	assign w325 = {w324, w323};
	assign w2849 = s305[31:31];
	assign w72 = {1'b0, w71};
	assign w2560 = w275 ? w2559 : w2558;
	assign w2850 = {w2849, w2848};
	assign w2851 = s305[31:31];
	assign w3082 = i13;
	assign w2853 = s305[31:31];
	assign w2855 = s305[31:31];
	assign w2858 = {w2857, w2856};
	assign w1403 = w1297[33:33];
	assign w1318 = w1245;
	assign w2861 = s305[31:31];

	// array write assignments
	always_comb begin
	end


	// state updates and reset
	always @(posedge clk) begin
		if (rst) begin
			s3047 <= w3046;
			s2626 <= w2625;
			s2601 <= w47;
			s2597 <= w117;
			s118 <= w117;
			s123 <= w47;
			s2700 <= w47;
			s1492 <= w791;
			s2606 <= w2605;
			s305 <= w304;
			s1043 <= w1042;
			s3040 <= w3039;
			s404 <= w403;
			s1007 <= w1006;
			s2618 <= w117;
			s772 <= w47;
			s792 <= w791;
			s797 <= w791;
			s409 <= w403;
			s1069 <= w1068;
			s1011 <= w1010;
		end
		else begin
			s3047 <= w4991;
			s3011 <= w4985;
			s3006 <= w4982;
			s3001 <= w4979;
			s2999 <= w4954;
			s2995 <= w4935;
			s2971 <= w4930;
			s2760 <= w4927;
			s2729 <= w4899;
			s2705 <= w4894;
			s2632 <= w4885;
			s2618 <= w4876;
			s2617 <= w4873;
			s2615 <= w4870;
			s2612 <= w4867;
			s2611 <= w4863;
			s2606 <= w4850;
			s2597 <= w4835;
			s2001 <= w4829;
			s2000 <= w4825;
			s1998 <= w4821;
			s1997 <= w4817;
			s1994 <= w4813;
			s1993 <= w4809;
			s1991 <= w4805;
			s1985 <= w4793;
			s1983 <= w4789;
			s1979 <= w4781;
			s1976 <= w4773;
			s1967 <= w4756;
			s1966 <= w4752;
			s1962 <= w4744;
			s1955 <= w4732;
			s1954 <= w4728;
			s1952 <= w4724;
			s1951 <= w4720;
			s1947 <= w4712;
			s1945 <= w4708;
			s1990 <= w4801;
			s1938 <= w4699;
			s1931 <= w4683;
			s1930 <= w4679;
			s1927 <= w4671;
			s1920 <= w4659;
			s1919 <= w4655;
			s1937 <= w4695;
			s1915 <= w4647;
			s1912 <= w4639;
			s1907 <= w4634;
			s1904 <= w4626;
			s1900 <= w4618;
			s1899 <= w4614;
			s1897 <= w4610;
			s1896 <= w4606;
			s1892 <= w4602;
			s1891 <= w4598;
			s1888 <= w4590;
			s1885 <= w4586;
			s1884 <= w4582;
			s1882 <= w4578;
			s1874 <= w4568;
			s1873 <= w4564;
			s1871 <= w4560;
			s1867 <= w4552;
			s1864 <= w4544;
			s1859 <= w4536;
			s1934 <= w4687;
			s1855 <= w4524;
			s1852 <= w4520;
			s1849 <= w4512;
			s1843 <= w4503;
			s1579 <= w3962;
			s1570 <= w3942;
			s1568 <= w3938;
			s1679 <= w4168;
			s1561 <= w3922;
			s1491 <= w3765;
			s1808 <= w4430;
			s1560 <= w3918;
			s439 <= w3365;
			s1546 <= w3895;
			s1467 <= w3721;
			s1537 <= w3875;
			s1735 <= w4282;
			s1534 <= w3867;
			s1528 <= w3855;
			s1521 <= w3844;
			s1660 <= w4128;
			s2991 <= w4933;
			s1764 <= w4337;
			s1796 <= w4406;
			s1542 <= w3883;
			s1520 <= w3839;
			s1514 <= w3823;
			s1839 <= w4491;
			s1923 <= w4667;
			s1513 <= w3818;
			s1975 <= w4769;
			s1632 <= w4067;
			s1571 <= w3946;
			s900 <= w3540;
			s1504 <= w3796;
			s2700 <= w4888;
			s468 <= w3428;
			s1744 <= w4302;
			s1916 <= w4651;
			s1866 <= w4548;
			s1501 <= w3786;
			s1578 <= w3958;
			s2626 <= w4881;
			s1575 <= w3950;
			s1719 <= w4246;
			s1497 <= w3779;
			s1490 <= w3758;
			s1305 <= w3715;
			s1270 <= w3678;
			s1647 <= w4099;
			s1773 <= w4357;
			s1535 <= w3871;
			s1201 <= w3624;
			s1550 <= w3903;
			s1682 <= w4176;
			s1191 <= w3622;
			s1160 <= w3618;
			s1127 <= w3574;
			s1069 <= w3572;
			s762 <= w3497;
			s885 <= w3525;
			s1518 <= w3834;
			s455 <= w3401;
			s1640 <= w4083;
			s1836 <= w4487;
			s960 <= w3546;
			s1595 <= w3996;
			s1007 <= w3554;
			s1527 <= w3851;
			s2601 <= w4842;
			s415 <= w3315;
			s1922 <= w4663;
			s896 <= w3529;
			s440 <= w3369;
			s437 <= w3357;
			s1134 <= w3582;
			s1549 <= w3899;
			s1635 <= w4075;
			s1517 <= w3829;
			s1234 <= w3666;
			s1913 <= w4643;
			s22 <= w3199;
			s475 <= w3457;
			s1948 <= w4716;
			s297 <= w3278;
			s1543 <= w3887;
			s1777 <= w4365;
			s416 <= w3321;
			s1616 <= w4040;
			s1828 <= w4471;
			s180 <= w3259;
			s458 <= w3414;
			s1840 <= w4495;
			s1944 <= w4704;
			s1553 <= w3911;
			s49 <= w3204;
			s235 <= w3266;
			s409 <= w3288;
			s1726 <= w4262;
			s31 <= w3202;
			s1856 <= w4528;
			s421 <= w3346;
			s118 <= w3224;
			s474 <= w3453;
			s1617 <= w4044;
			s404 <= w3284;
			s2609 <= w4859;
			s441 <= w3374;
			s1982 <= w4785;
			s1745 <= w4306;
			s453 <= w3393;
			s772 <= w3504;
			s109 <= w3220;
			s1207 <= w3631;
			s420 <= w3342;
			s1698 <= w4205;
			s55 <= w3216;
			s1848 <= w4508;
			s1663 <= w4132;
			s417 <= w3327;
			s107 <= w3218;
			s1928 <= w4675;
			s1858 <= w4532;
			s1530 <= w3859;
			s1538 <= w3879;
			s1254 <= w3669;
			s1710 <= w4229;
			s470 <= w3436;
			s1614 <= w4036;
			s1505 <= w3801;
			s471 <= w3440;
			s1641 <= w4087;
			s1889 <= w4594;
			s1043 <= w3567;
			s19 <= w2957;
			s1707 <= w4225;
			s418 <= w3332;
			s1960 <= w4740;
			s1729 <= w4270;
			s1795 <= w4402;
			s438 <= w3361;
			s1741 <= w4294;
			s1511 <= w3813;
			s1613 <= w4032;
			s2997 <= w4945;
			s1780 <= w4373;
			s152 <= w3246;
			s1656 <= w4116;
			s121 <= w3231;
			s469 <= w3432;
			s769 <= w3499;
			s2600 <= w4839;
			s984 <= w3550;
			s1650 <= w4107;
			s792 <= w3508;
			s1545 <= w3891;
			s1563 <= w3926;
			s1792 <= w4394;
			s419 <= w3338;
			s1758 <= w4325;
			s1552 <= w3907;
			s305 <= w3280;
			s18 <= w3172;
			s457 <= w3410;
			s2702 <= w4891;
			s127 <= w736;
			s813 <= w3518;
			s1625 <= w4051;
			s1531 <= w3863;
			s443 <= w3382;
			s1609 <= w4024;
			s1935 <= w4691;
			s1294 <= w3712;
			s1703 <= w4213;
			s1789 <= w4390;
			s1502 <= w3791;
			s444 <= w3386;
			s898 <= w3531;
			s815 <= w3521;
			s456 <= w3405;
			s459 <= w3418;
			s1842 <= w4499;
			s473 <= w3449;
			s1659 <= w4124;
			s1881 <= w4574;
			s1870 <= w4556;
			s1738 <= w4290;
			s1628 <= w4059;
			s1582 <= w3966;
			s1755 <= w4317;
			s1835 <= w4483;
			s1827 <= w4467;
			s1583 <= w3970;
			s1626 <= w4055;
			s1754 <= w4313;
			s1633 <= w4071;
			s1585 <= w3974;
			s1592 <= w3988;
			s1594 <= w3992;
			s1598 <= w4000;
			s1903 <= w4622;
			s1599 <= w4004;
			s1959 <= w4736;
			s1821 <= w4455;
			s1601 <= w4008;
			s1978 <= w4777;
			s1576 <= w3954;
			s797 <= w3514;
			s1678 <= w4164;
			s1602 <= w4012;
			s1606 <= w4016;
			s1607 <= w4020;
			s1610 <= w4028;
			s1851 <= w4516;
			s1586 <= w3978;
			s1629 <= w4063;
			s1636 <= w4079;
			s1492 <= w3514;
			s1643 <= w4091;
			s1762 <= w4333;
			s1644 <= w4095;
			s1648 <= w4103;
			s1651 <= w4111;
			s1863 <= w4540;
			s1657 <= w4120;
			s1671 <= w4148;
			s1970 <= w4764;
			s1672 <= w4152;
			s1675 <= w4160;
			s1681 <= w4172;
			s1906 <= w4630;
			s1688 <= w4181;
			s1691 <= w4189;
			s1674 <= w4156;
			s1692 <= w4193;
			s3000 <= w4970;
			s442 <= w3378;
			s1737 <= w4286;
			s239 <= w3268;
			s1742 <= w4298;
			s1695 <= w4197;
			s3040 <= w4988;
			s1696 <= w4201;
			s1699 <= w4209;
			s1704 <= w4217;
			s1264 <= w3671;
			s1714 <= w4241;
			s1706 <= w4221;
			s1667 <= w4144;
			s1711 <= w4233;
			s1713 <= w4237;
			s1496 <= w3773;
			s1720 <= w4250;
			s422 <= w3350;
			s1689 <= w4185;
			s1722 <= w4254;
			s1730 <= w4274;
			s123 <= w3234;
			s1820 <= w4451;
			s1723 <= w4258;
			s1727 <= w4266;
			s1963 <= w4748;
			s1734 <= w4278;
			s1969 <= w4760;
			s1757 <= w4321;
			s1761 <= w4329;
			s1765 <= w4341;
			s1664 <= w4136;
			s454 <= w3397;
			s1769 <= w4345;
			s1770 <= w4349;
			s1772 <= w4353;
			s1510 <= w3808;
			s1776 <= w4361;
			s1779 <= w4369;
			s1785 <= w4378;
			s1567 <= w3934;
			s1786 <= w4382;
			s1986 <= w4797;
			s1788 <= w4386;
			s1810 <= w4434;
			s1793 <= w4398;
			s1800 <= w4410;
			s460 <= w3422;
			s1801 <= w4414;
			s1564 <= w3930;
			s1803 <= w4418;
			s1666 <= w4140;
			s1804 <= w4422;
			s472 <= w3445;
			s1807 <= w4426;
			s1811 <= w4438;
			s1817 <= w4443;
			s1818 <= w4447;
			s1824 <= w4459;
			s2596 <= w4832;
			s1591 <= w3984;
			s1825 <= w4463;
			s1011 <= w3559;
			s1832 <= w4475;
			s1833 <= w4479;
		end
	end

	// assumptions
	always @* begin
		assume (w533);
		assume (w682);
		assume (w685);
	end;

	// assertions
	always @* begin
		assert (~w542);
	end
endmodule


