`timescale 1ns / 1ps

/*
mriscvcore
by CKDUR

This is the definitive core.
*/
module top(
   input clk,
   input [31:0] instruction,
   input rstn,
   input outside_resetn,
    input [31:0] Rdata,
    input ARready,
    input Rvalid,
    input AWready,
    input Wready,
    input Bvalid, 
    output [31:0] AWdata,
    output [31:0] ARdata,
    output [31:0] Wdata,
    output ARvalid,
    output RReady,
    output AWvalid,
    output Wvalid,
    output [2:0] ARprot,AWprot,
    output Bready,
    output [3:0] Wstrb,
    
    // IRQ interface
    
    input [31:0] inirr,
    output [31:0] outirr,
    output trap
);
   inst_constraint inst_constraint0(.clk(clk),
                                    .instruction(instruction));
	always @* begin
		no_reset: assume(outside_resetn);
	end
   assume property (Rdata==32'b0);
   mriscvcore RTL(
    .clk(clk),
    .instruction(instruction),
    .rstn(rstn),
    .outside_resetn(outside_resetn),
    .Rdata(Rdata),
    .ARready(ARready),
    .Rvalid(Rvalid),
    .AWready(AWready),
    .Wready(Wready),
    .Bvalid(Bvalid),
    .AWdata(AWdata),
    .ARdata(ARdata),
    .Wdata(Wdata),
    .ARvalid(ARvalid),
    .RReady(RReady),
    .AWvalid(AWvalid),
    .Wvalid(Wvalid),
    .ARprot(ARprot),
    .AWprot(AWprot),
    .Bready(Bready),
    .Wstrb(Wstrb),
    .inirr(inirr),
    .outirr(outirr),
    .trap(trap)
   );
endmodule



module mriscvcore(
    input clk,
    input [31:0] instruction,
    input rstn,
    input outside_resetn,
    // AXI-4 LITE INTERFACE
    input [31:0] Rdata,
    input ARready,
    input Rvalid,
    input AWready,
    input Wready,
    input Bvalid, 
    output [31:0] AWdata,
    output [31:0] ARdata,
    output [31:0] Wdata,
    output ARvalid,
    output RReady,
    output AWvalid,
    output Wvalid,
    output [2:0] ARprot,AWprot,
    output Bready,
    output [3:0] Wstrb,
    
    // IRQ interface
    
    input [31:0] inirr,
    output [31:0] outirr,
    output trap
     
    );
    
// SIGNAL DECLARATION     *********************************************************

// Data Buses
wire [31:0] rd, rs1, rs2, imm, pc, inst, qed_ifu_instruction;
wire [11:0] code;
wire [11:0] codif;

// Auxiliars
wire [4:0] rs1i, rs2i, rdi;

//IRQ SIGNALS
wire [31:0] pc_c, addrm, pc_irq;
wire flag;
//MEMORY INTERFACE SIGNALS
wire is_rd_mem;
wire [1:0] W_R_mem, wordsize_mem;
wire sign_mem, en_mem, busy_mem, done_mem, align_mem;
//SIGNALS DECO INST
wire enableDec;    
//SIGNALS MULT
wire enable_mul, done_mul, is_inst_mul;
//SIGNALS ALU
wire cmp, carry, enable_alu, is_inst_alu, is_rd_alu;
//SIGNALS UTILITY
wire is_inst_util, is_rd_util;
//SIGNALS FSM
wire is_exec;
wire qed_vld_out;
wire qed_vld_out_q;

// DATAPATH PHASE    *************************************************************

MEMORY_INTERFACE MEMORY_INTERFACE_inst(
    .clock(clk),
    .resetn(rstn),
    .outside_resetn(outside_resetn),
    .instruction(instruction),
    .rdw_rsrn(rdw_rsrn),
    // Data buses
    .rs1(rs1),
    .rs2(rs2),
    .rd(rd),
    .imm(imm), 
    .pc(pc),
    .rd_en(is_rd_mem),
    // AXI4-Interface
    .Rdata_mem(Rdata),
    .ARready(ARready),
    .Rvalid(Rvalid),
    .AWready(AWready),
    .Wready(Wready),
    .Bvalid(Bvalid),
    .AWdata(AWdata),
    .ARdata(ARdata),
    .Wdata(Wdata),
    .ARvalid(ARvalid),
    .RReady(RReady),
    .AWvalid(AWvalid),
    .Wvalid(Wvalid),
    .arprot(ARprot),
    .awprot(AWprot),
    .Bready(Bready),
    .Wstrb(Wstrb),
    // To DECO_INSTR
    .inst(inst),
    .qed_ifu_instruction_o(qed_ifu_instruction),
    // To FSM
    .W_R(W_R_mem),
    .wordsize(wordsize_mem),
    .signo(sign_mem),
    .enable(en_mem),
    .busy(busy_mem), 
    .done(done_mem),
    .align(align_mem),
    .qed_vld_out(qed_vld_out)
    );


DECO_INSTR DECO_INSTR_inst(
    .clk(clk),
    // From MEMORY_INTERFACE
    .inst(qed_ifu_instruction),
    // Auxiliars to BUS
    .rs1i(rs1i),
    .rs2i(rs2i),
    .rdi(rdi),
    .imm(imm),
    .code(code),
    .codif(codif)
    );

REG_FILE REG_FILE_inst(
    .clk(clk),
    .rst(rstn),
    .outside_resetn(outside_resetn),
    .qed_vld_out_q(qed_vld_out_q),
    .rd(rd),
    .rdi(rdi),
    .rdw_rsrn(rdw_rsrn),
    .rs1(rs1),
    .rs1i(rs1i),
    .rs2(rs2),
    .rs2i(rs2i)
    );

    
ALU ALU_inst(
    .clk(clk),
    .reset(rstn),
    // Data Buses
    .rs1(rs1),
    .rs2(rs2),
    .rd(rd),
    .decinst(code),
    .imm(imm),
    // To UTILITY
    .cmp(cmp),
    // To FSM
    .en(enable_alu),
    .carry(carry),
    .is_rd(is_rd_alu),
    .is_inst(is_inst_alu)
    );
    
     
IRQ IRQ_inst(
    .rst(rstn),
    .clk(clk),
    .savepc(1'b0),
    .en(1'b0),
    .instr(code),
    .rs1(rs1),
    .rs2(rs2),
    .inirr(inirr),
    .pc(pc),
    .imm(imm),
    .rd(rd),
    .addrm(addrm),
    .outirr(outirr),
    .pc_irq(pc_irq),
    .pc_c(pc_c),
    .flag(flag)
    );

MULT MULT_inst(
    .clk(clk),
    .reset(rstn),
    .rs1(rs1),
    .rs2(rs2),
    .rd(rd),
    .Enable(enable_mul),
    .is_oper(is_inst_mul),
    .Done(done_mul),
    .codif(code)
    );

UTILITY UTILITY_inst(
    .clk(clk),
    .rst(rstn),
    // FROM DATA BUS
    .rs1(rs1),
    .rd(rd),
    .opcode(code),
    .imm(imm),
    .pc(pc),
    // FROM IRQ
    .irr_ret(pc_c),
    .irr_dest(pc_irq),
    // FROM ALU
    .branch(cmp),
    // FSM
    .irr(1'b0),
    .enable_pc(enable_pc),
    .is_inst(is_inst_util),
    .is_rd(is_rd_util)
    );

// FINITE-STATE MACHINE PHASE    *************************************************

FSM FSM_inst
    (
    .clk(clk),
    .reset(rstn),
    .outside_resetn(outside_resetn),
    .qed_vld_out(qed_vld_out),
    // Auxiliars from DATAPATH
    .codif(codif),
    
    // Inputs from DATAPATH
    .busy_mem(busy_mem), 
    .done_mem(done_mem),
    .aligned_mem(align_mem),
    .done_exec(done_exec),
    .is_exec(is_exec),
    
    // Outputs to DATAPATH
    .W_R_mem(W_R_mem),
    .wordsize_mem(wordsize_mem),
    .sign_mem(sign_mem),
    .en_mem(en_mem),
    .enable_exec(enable_exec),
    .enable_exec_mem(enable_exec_mem),
    .trap(trap),
    .enable_pc(enable_pc),
    .qed_vld_out_q(qed_vld_out_q)
    );
    
    // Enable Assign
    assign enable_mul = enable_exec; 
    assign enable_alu = enable_exec;
    
    // Done Assign
    assign done_exec = is_inst_util | is_inst_alu | (done_mul & is_inst_mul);
    
    // Is exec assign
    assign is_exec = ~(&(code));
    
    // Write to rd flag
    assign rdw_rsrn = (is_rd_util | is_rd_alu | done_mul | (is_rd_mem & done_mem)) & (enable_exec | enable_exec_mem);

endmodule

